* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
*.PININFO A1:I A2:I Z:O VDD:P VNW:P VPW:P VSS:G
*.EQN Z=!((A1 * A2) + !(A1 + A2))
M_i_6 I A2 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_7 VSS A1 I VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_2 Z I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 net_0 A1 Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8 net_2 A2 I VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_9 VDD A1 net_2 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_5 net_1 I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3 Z A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4 net_1 A2 Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
