# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.3 1.77 9.93 1.77 9.93 2.27 11.23 2.27 11.23 2.5 9.3 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.75 2.215 0.98 2.215 0.98 2.73 3.51 2.73 3.51 2.27 4.13 2.27 4.13 2.73 8.125 2.73 8.125 2.215 8.355 2.215 8.355 2.96 0.75 2.96  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 1.81 4.64 1.81 4.64 2.27 6.27 2.27 6.27 2.5 4.41 2.5 4.41 2.04 1.99 2.04 1.99 2.5 1.21 2.5  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.22 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 3.19 11.965 3.19 11.965 1.515 9.825 1.515 9.825 1.14 10.055 1.14 10.055 1.285 12.01 1.285 12.01 1.14 12.79 1.14 12.79 1.53 12.195 1.53 12.195 4.36 11.965 4.36 11.965 3.42 9.955 3.42 9.955 4.36 9.725 4.36 9.725 3.42 7.915 3.42 7.915 4.36 7.685 4.36 7.685 3.42 5.775 3.42 5.775 4.36 5.545 4.36 5.545 3.42 3.635 3.42 3.635 4.36 3.405 4.36 3.405 3.42 1.495 3.42 1.495 4.36 1.265 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.65 0.475 3.65 0.475 4.59 2.285 4.59 2.285 3.875 2.515 3.875 2.515 4.59 4.425 4.59 4.425 3.65 4.655 3.65 4.655 4.59 6.565 4.59 6.565 3.65 6.795 3.65 6.795 4.59 8.705 4.59 8.705 3.65 8.935 3.65 8.935 4.59 10.845 4.59 10.845 3.65 11.075 3.65 11.075 4.59 13.085 4.59 13.085 3.65 13.315 3.65 13.315 4.59 13.415 4.59 14 4.59 14 5.49 13.415 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14 -0.45 14 0.45 6.895 0.45 6.895 1.11 6.665 1.11 6.665 0.45 2.615 0.45 2.615 1.11 2.385 1.11 2.385 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.77 0.475 0.77 0.475 1.35 2.845 1.35 2.845 0.77 4.755 0.77 4.755 1.35 8.94 1.35 8.94 0.68 13.415 0.68 13.415 1.58 13.185 1.58 13.185 0.91 11.23 0.91 11.23 1.055 10.89 1.055 10.89 0.91 9.17 0.91 9.17 1.58 4.525 1.58 4.525 1 3.075 1 3.075 1.58 0.245 1.58  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nand3_4
