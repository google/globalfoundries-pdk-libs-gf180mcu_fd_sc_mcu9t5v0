# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.84 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 2.33 3.895 2.33 3.895 2.71 2.945 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.105 1.21 14.41 1.21 14.41 1.59 14.335 1.59 14.335 2.05 14.105 2.05  ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.235 1.575 2.235 1.575 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.685 2.875 19.485 2.875 19.715 2.875 19.715 1.655 17.685 1.655 17.685 0.845 17.915 0.845 17.915 1.395 19.75 1.395 19.75 0.815 20.175 0.815 20.175 3.685 19.725 3.685 19.725 3.295 19.485 3.295 17.915 3.295 17.915 3.685 17.685 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.225 4.59 3.225 3.615 3.455 3.615 3.455 4.59 5.99 4.59 7.305 4.59 7.305 3.615 7.535 3.615 7.535 4.59 8.555 4.59 9.045 4.59 9.045 3.38 9.275 3.38 9.275 4.59 9.77 4.59 10.295 4.59 13.525 4.59 13.525 4.345 13.755 4.345 13.755 4.59 15.55 4.59 15.845 4.59 15.845 3.875 16.075 3.875 16.075 4.59 16.665 4.59 16.665 3.875 16.895 3.875 16.895 4.59 18.705 4.59 18.705 3.875 18.935 3.875 18.935 4.59 19.485 4.59 20.745 4.59 20.745 3.875 20.975 3.875 20.975 4.59 21.84 4.59 21.84 5.49 19.485 5.49 15.55 5.49 10.295 5.49 9.77 5.49 8.555 5.49 5.99 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.84 -0.45 21.84 0.45 21.275 0.45 21.275 1.165 21.045 1.165 21.045 0.45 19.035 0.45 19.035 1.165 18.805 1.165 18.805 0.45 16.795 0.45 16.795 1.165 16.565 1.165 16.565 0.45 13.655 0.45 13.655 1.25 13.425 1.25 13.425 0.45 8.955 0.45 8.955 1.25 8.725 1.25 8.725 0.45 3.435 0.45 3.435 1.25 3.205 1.25 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.245 1.25 4.555 1.25 4.555 3.785 4.245 3.785  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 3.155 3.915 3.155 3.915 4.13 5.99 4.13 5.99 4.36 3.685 4.36 3.685 3.385 2.615 3.385 2.615 3.685 2.385 3.685  ;
        POLYGON 6.285 3.145 8.555 3.145 8.555 3.955 8.325 3.955 8.325 3.375 6.515 3.375 6.515 3.955 6.285 3.955  ;
        POLYGON 5.265 1.25 5.675 1.25 5.675 2.685 9.77 2.685 9.77 2.915 5.495 2.915 5.495 3.785 5.265 3.785  ;
        POLYGON 6.81 2.225 10.065 2.225 10.065 1.25 10.295 1.25 10.295 4.02 10.065 4.02 10.065 2.455 6.81 2.455  ;
        POLYGON 6.07 1.765 9.605 1.765 9.605 0.79 11.875 0.79 11.875 3.09 11.645 3.09 11.645 1.02 10.755 1.02 10.755 2.05 10.525 2.05 10.525 1.02 9.835 1.02 9.835 1.995 6.07 1.995  ;
        POLYGON 12.285 1.25 12.535 1.25 12.535 3.55 12.285 3.55  ;
        POLYGON 11.185 1.25 11.415 1.25 11.415 3.21 11.42 3.21 11.42 3.79 15.07 3.79 15.07 2.47 15.55 2.47 15.55 2.7 15.3 2.7 15.3 4.02 11.185 4.02  ;
        POLYGON 12.81 2.32 14.61 2.32 14.61 2.01 15.845 2.01 15.845 0.845 16.075 0.845 16.075 2.015 19.485 2.015 19.485 2.275 15.845 2.275 15.845 2.24 14.84 2.24 14.84 3.215 14.555 3.215 14.555 2.55 12.81 2.55  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4
