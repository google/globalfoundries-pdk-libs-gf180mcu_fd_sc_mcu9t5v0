* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__icgtn_4 CLKN E TE Q VDD VNW VPW VSS
*.PININFO CLKN:I E:I TE:I Q:O VDD:P VNW:P VPW:P VSS:G
M_MU19 VSS TE net50 VPW nfet_05v0 W=0.700000U L=0.600000U
M_MU20 net50 E VSS VPW nfet_05v0 W=0.700000U L=0.600000U
M_MI82 net53 NCP net50 VPW nfet_05v0 W=0.700000U L=0.600000U
M_MI91 net038 CP net53 VPW nfet_05v0 W=0.700000U L=0.600000U
M_MI92 VSS QD net038 VPW nfet_05v0 W=0.700000U L=0.600000U
M_MU82_M_u2 NCP CP VSS VPW nfet_05v0 W=0.700000U L=0.600000U
M_MI95_M_u2 VSS net53 QD VPW nfet_05v0 W=0.700000U L=0.600000U
M_MI89_M_u2 net36 QD VSS VPW nfet_05v0 W=0.700000U L=0.600000U
M_MU81_M_u2 VSS CLKN CP VPW nfet_05v0 W=0.800000U L=0.600000U
M_MI1_M_u3 d3 net36 VSS VPW nfet_05v0 W=0.800000U L=0.600000U
M_MI1_M_u4 VSS CLKN d3 VPW nfet_05v0 W=0.800000U L=0.600000U
M_MU75_M_u2 Q d3 VSS VPW nfet_05v0 W=1.000000U L=0.600000U
M_MU75_M_u2_19 Q d3 VSS VPW nfet_05v0 W=1.000000U L=0.600000U
M_MU75_M_u2_33 Q d3 VSS VPW nfet_05v0 W=1.000000U L=0.600000U
M_MU75_M_u2_19_5 Q d3 VSS VPW nfet_05v0 W=1.000000U L=0.600000U
M_MI81 net58 TE VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_MU17 net61 E net58 VNW pfet_05v0 W=1.380000U L=0.500000U
M_MU16 net53 CP net61 VNW pfet_05v0 W=1.380000U L=0.500000U
M_MI90 net067 NCP net53 VNW pfet_05v0 W=1.380000U L=0.500000U
M_MI88 VDD QD net067 VNW pfet_05v0 W=1.380000U L=0.500000U
M_MU82_M_u3 NCP CP VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_MI95_M_u3 VDD net53 QD VNW pfet_05v0 W=1.380000U L=0.500000U
M_MI89_M_u3 net36 QD VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_MU81_M_u3 VDD CLKN CP VNW pfet_05v0 W=1.680000U L=0.500000U
M_MI1_M_u1 XI1-net8 net36 VDD VNW pfet_05v0 W=1.680000U L=0.500000U
M_MI1_M_u2 d3 CLKN XI1-net8 VNW pfet_05v0 W=1.680000U L=0.500000U
M_MU75_M_u3 Q d3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_MU75_M_u3_1 Q d3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_MU75_M_u3_2 Q d3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_MU75_M_u3_1_35 Q d3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
