* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__addh_2 A B CO S VDD VNW VPW VSS
*.PININFO A:I B:I CO:O S:O VDD:P VNW:P VPW:P VSS:G
*.EQN CO=(A * B);S=!((A * B) + !(A + B))
M_i_2_1 CO NCO VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 VSS NCO CO VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5 net_0 A VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4 NCO B net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9 NS B net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8 net_1 A NS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10 VSS NCO net_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 S NS VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 VSS NS S VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 CO NCO VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 VDD NCO CO VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7 NCO A VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 VDD B NCO VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_12 net_2 B VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11 NS A net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_13 VDD NCO NS VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 S NS VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 VDD NS S VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
