# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 29.12 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.076 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.57 1.785 6.01 1.785 6.01 3.27 5.57 3.27  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.2744 ;
    PORT
      LAYER METAL1 ;
        POLYGON 16.14 3.01 25.57 3.01 25.94 3.01 26.45 3.01 26.45 1.595 16.09 1.595 16.09 0.895 27.52 0.895 27.52 1.595 26.98 1.595 26.98 3.01 26.97 3.01 26.97 4.28 26.735 4.28 26.735 3.49 25.94 3.49 25.57 3.49 24.93 3.49 24.93 4.28 24.7 4.28 24.7 3.49 22.89 3.49 22.89 4.28 22.66 4.28 22.66 3.49 20.75 3.49 20.75 4.28 20.52 4.28 20.52 3.49 18.51 3.49 18.51 4.28 18.28 4.28 18.28 3.49 16.37 3.49 16.37 4.28 16.14 4.28  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.83 4.59 1.83 3.47 2.06 3.47 2.06 4.59 6.03 4.59 6.03 4.51 6.26 4.51 6.26 4.59 8.51 4.59 8.51 4.51 8.74 4.51 8.74 4.59 10.77 4.59 10.77 3.95 11 3.95 11 4.59 12.81 4.59 12.81 3.47 13.04 3.47 13.04 4.59 14.92 4.59 14.92 3.88 15.15 3.88 15.15 4.59 17.16 4.59 17.16 3.96 17.39 3.96 17.39 4.59 19.4 4.59 19.4 3.94 19.63 3.94 19.63 4.59 21.64 4.59 21.64 3.94 21.87 3.94 21.87 4.59 23.68 4.59 23.68 3.94 23.91 3.94 23.91 4.59 25.57 4.59 25.72 4.59 25.72 3.94 25.94 3.94 25.95 3.94 25.95 4.59 27.76 4.59 27.76 3.47 27.99 3.47 27.99 4.59 29.12 4.59 29.12 5.49 25.94 5.49 25.57 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 29.12 -0.45 29.12 0.45 28.64 0.45 28.64 1.54 28.41 1.54 28.41 0.45 26.455 0.45 26.455 0.635 26.115 0.635 26.115 0.45 24.215 0.45 24.215 0.635 23.875 0.635 23.875 0.45 21.975 0.45 21.975 0.635 21.635 0.635 21.635 0.45 19.735 0.45 19.735 0.635 19.395 0.635 19.395 0.45 17.495 0.45 17.495 0.635 17.155 0.635 17.155 0.45 15.2 0.45 15.2 1.54 14.97 1.54 14.97 0.45 12.96 0.45 12.96 1.54 12.73 1.54 12.73 0.45 10.72 0.45 10.72 1.54 10.49 1.54 10.49 0.45 8.535 0.45 8.535 0.635 8.195 0.635 8.195 0.45 6.295 0.45 6.295 0.635 5.955 0.635 5.955 0.45 1.595 0.45 1.595 1.07 1.365 1.07 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.81 2.94 1.805 2.94 1.805 1.54 0.245 1.54 0.245 0.73 0.475 0.73 0.475 1.31 2.035 1.31 2.035 2.48 3.575 2.48 3.575 3.17 1.04 3.17 1.04 4.28 0.81 4.28  ;
        POLYGON 4.79 3.01 5.02 3.01 5.02 3.59 7.27 3.59 7.27 2.23 8.69 2.23 8.69 1.555 4.835 1.555 4.835 1.325 8.975 1.325 8.975 2.525 7.5 2.525 7.5 3.82 4.79 3.82  ;
        POLYGON 2.85 3.47 3.08 3.47 3.08 4.05 4.33 4.05 4.33 1.595 3.55 1.595 3.55 1.365 4.56 1.365 4.56 4.05 9.75 4.05 9.75 2.505 25.57 2.505 25.57 2.735 14.06 2.735 14.06 4.28 13.83 4.28 13.83 2.735 12.02 2.735 12.02 4.28 11.79 4.28 11.79 2.735 9.98 2.735 9.98 4.28 2.85 4.28  ;
        POLYGON 2.485 0.73 2.715 0.73 2.715 0.865 9.315 0.865 9.315 0.815 9.66 0.815 9.66 1.825 11.61 1.825 11.61 0.84 11.84 0.84 11.84 1.825 13.85 1.825 13.85 0.84 14.08 0.84 14.08 1.825 25.94 1.825 25.94 2.055 9.43 2.055 9.43 1.095 3.32 1.095 3.32 1.825 4.1 1.825 4.1 3.82 3.87 3.82 3.87 2.055 3.09 2.055 3.09 1.095 2.715 1.095 2.715 1.54 2.485 1.54  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_12
