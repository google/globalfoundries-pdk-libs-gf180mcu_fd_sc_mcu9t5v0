# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.135 1.77 2.135 2.555 1.83 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 1.77 3.26 1.77 3.26 2.5 2.92 2.5  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.99 1.77 4.33 1.77 4.33 2.5 3.99 2.5  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.6145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.77 0.97 1.77 0.97 2.5 0.63 2.5  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.5256 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.465 3.45 2.42 3.45 2.42 1.14 2.77 1.14 2.77 1.31 3.835 1.31 4.725 1.31 4.725 0.73 4.955 0.73 4.955 1.54 3.835 1.54 2.65 1.54 2.65 3.83 1.695 3.83 1.695 4.36 1.465 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 3.835 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 5.6 4.59 5.6 5.49 3.835 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 0.475 0.45 0.475 1.54 0.245 1.54 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 0.68 3.835 0.68 3.835 1.07 3.605 1.07 3.605 0.91 1.595 0.91 1.595 1.54 1.365 1.54  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_1
