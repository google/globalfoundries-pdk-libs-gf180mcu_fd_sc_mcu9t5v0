# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 36.96 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.815 1.85 1.155 1.85 1.155 2.275 0.815 2.275  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.768 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.065 2.03 7.71 2.03 7.71 2.605 5.065 2.605  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 14.3292 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.405 2.965 33.7 2.965 33.73 2.965 34.835 2.965 34.835 1.595 19.405 1.595 19.405 0.895 35.315 0.895 35.315 4.12 35.085 4.12 35.085 3.365 33.73 3.365 33.7 3.365 32.975 3.365 32.975 4.12 32.745 4.12 32.745 3.365 30.735 3.365 30.735 4.12 30.505 4.12 30.505 3.365 28.495 3.365 28.495 4.12 28.265 4.12 28.265 3.365 26.255 3.365 26.255 4.12 26.025 4.12 26.025 3.365 24.015 3.365 24.015 4.12 23.785 4.12 23.785 3.365 21.775 3.365 21.775 4.12 21.545 4.12 21.545 3.365 19.635 3.365 19.635 4.12 19.405 4.12  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.905 4.59 1.905 3.31 2.135 3.31 2.135 4.59 4.665 4.59 4.665 4.35 4.895 4.35 4.895 4.59 6.805 4.59 6.805 4.35 7.035 4.35 7.035 4.59 9.045 4.59 9.045 3.31 9.275 3.31 9.275 4.59 11.285 4.59 11.285 3.31 11.515 3.31 11.515 4.59 13.525 4.59 13.525 3.31 13.755 3.31 13.755 4.59 15.765 4.59 15.765 3.31 15.995 3.31 15.995 4.59 18.185 4.59 18.185 3.88 18.415 3.88 18.415 4.59 20.425 4.59 20.425 3.745 20.655 3.745 20.655 4.59 22.665 4.59 22.665 3.745 22.895 3.745 22.895 4.59 24.905 4.59 24.905 3.745 25.135 3.745 25.135 4.59 27.145 4.59 27.145 3.745 27.375 3.745 27.375 4.59 29.385 4.59 29.385 3.745 29.615 3.745 29.615 4.59 31.625 4.59 31.625 3.745 31.855 3.745 31.855 4.59 33.7 4.59 33.73 4.59 33.865 4.59 33.865 3.745 34.095 3.745 34.095 4.59 36.105 4.59 36.105 3.31 36.335 3.31 36.335 4.59 36.96 4.59 36.96 5.49 33.73 5.49 33.7 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 36.96 -0.45 36.96 0.45 36.435 0.45 36.435 1.49 36.205 1.49 36.205 0.45 34.25 0.45 34.25 0.665 33.91 0.665 33.91 0.45 32.01 0.45 32.01 0.665 31.67 0.665 31.67 0.45 29.77 0.45 29.77 0.665 29.43 0.665 29.43 0.45 27.53 0.45 27.53 0.665 27.19 0.665 27.19 0.45 25.29 0.45 25.29 0.665 24.95 0.665 24.95 0.45 23.05 0.45 23.05 0.665 22.71 0.665 22.71 0.45 20.81 0.45 20.81 0.665 20.47 0.665 20.47 0.45 18.515 0.45 18.515 1.49 18.285 1.49 18.285 0.45 16.095 0.45 16.095 1.49 15.865 1.49 15.865 0.45 13.855 0.45 13.855 1.49 13.625 1.49 13.625 0.45 11.615 0.45 11.615 1.455 11.385 1.455 11.385 0.45 9.43 0.45 9.43 0.64 9.09 0.64 9.09 0.45 7.19 0.45 7.19 0.64 6.85 0.64 6.85 0.45 4.95 0.45 4.95 0.64 4.61 0.64 4.61 0.45 1.595 0.45 1.595 1.16 1.365 1.16 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.885 2.505 1.805 2.505 1.805 1.62 0.245 1.62 0.245 0.68 0.475 0.68 0.475 1.39 2.035 1.39 2.035 2.505 3.65 2.505 3.65 2.735 1.115 2.735 1.115 4.12 0.885 4.12  ;
        POLYGON 5.73 3.31 8.08 3.31 8.08 1.6 5.73 1.6 5.73 1.37 8.31 1.37 8.31 2.305 16.45 2.305 16.45 2.62 8.31 2.62 8.31 3.65 5.73 3.65  ;
        POLYGON 2.925 3.31 3.155 3.31 3.155 3.89 4.405 3.89 4.405 1.595 3.55 1.595 3.55 1.365 4.635 1.365 4.635 3.89 8.585 3.89 8.585 2.85 17.065 2.85 17.065 2.505 33.7 2.505 33.7 2.735 17.295 2.735 17.295 4.12 17.065 4.12 17.065 3.08 14.875 3.08 14.875 4.12 14.645 4.12 14.645 3.08 12.635 3.08 12.635 4.12 12.405 4.12 12.405 3.08 10.395 3.08 10.395 4.12 10.165 4.12 10.165 3.08 8.815 3.08 8.815 4.12 2.925 4.12  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.905 10.265 0.905 10.265 0.68 10.5 0.68 10.5 1.75 12.505 1.75 12.505 0.68 12.735 0.68 12.735 1.75 14.745 1.75 14.745 0.68 14.975 0.68 14.975 1.75 17.165 1.75 17.165 0.68 17.395 0.68 17.395 1.75 18.8 1.75 18.8 1.865 33.73 1.865 33.73 2.095 18.61 2.095 18.61 2.075 10.27 2.075 10.27 1.135 3.32 1.135 3.32 1.865 4.175 1.865 4.175 3.65 3.945 3.65 3.945 2.095 3.09 2.095 3.09 1.49 2.485 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_16
