# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 2.33 3.975 2.33 3.975 2.71 2.945 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.965 2.2 17.77 2.2 17.77 2.76 16.965 2.76  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.545 2.33 15.575 2.33 15.575 2.805 14.545 2.805  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.235 1.575 2.235 1.575 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.685 0.845 20.01 0.845 20.01 3.685 19.705 3.685 19.705 1.655 19.685 1.655  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.305 4.59 3.305 3.515 3.535 3.515 3.535 4.59 7.605 4.59 7.605 4.375 7.835 4.375 7.835 4.59 10.805 4.59 10.805 4.375 11.035 4.375 11.035 4.59 12.715 4.59 14.85 4.59 14.85 3.95 15.19 3.95 15.19 4.59 16.89 4.59 16.89 3.95 17.23 3.95 17.23 4.59 18.69 4.59 18.985 4.59 18.985 3.425 19.215 3.425 19.215 4.59 19.475 4.59 20.725 4.59 20.725 3.875 20.955 3.875 20.955 4.59 21.28 4.59 21.28 5.49 19.475 5.49 18.69 5.49 12.715 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 21.035 0.45 21.035 1.165 20.805 1.165 20.805 0.45 17.175 0.45 17.175 1.225 16.945 1.225 16.945 0.45 9.175 0.45 9.175 1.425 8.945 1.425 8.945 0.45 3.435 0.45 3.435 1.425 3.205 1.425 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 1.74 0.245 1.74 0.245 1.315 0.655 1.315 0.655 1.51 2.035 1.51 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.325 1.315 4.555 1.315 4.555 3.685 4.325 3.685  ;
        POLYGON 6.365 3.345 9.075 3.345 9.075 3.685 6.365 3.685  ;
        POLYGON 5.345 2.685 5.825 2.685 5.825 1.315 6.055 1.315 6.055 2.685 10.005 2.685 10.005 2.575 10.235 2.575 10.235 2.915 5.575 2.915 5.575 3.685 5.345 3.685  ;
        POLYGON 9.565 3.345 11.39 3.345 11.39 2.345 7.335 2.345 7.335 2.455 7.105 2.455 7.105 2.115 11.425 2.115 11.425 1.315 11.655 1.315 11.655 3.445 12.045 3.445 12.045 2.875 12.275 2.875 12.275 3.685 9.565 3.685  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 3.055 3.995 3.055 3.995 3.915 12.715 3.915 12.715 4.315 12.485 4.315 12.485 4.145 6.07 4.145 6.07 4.26 3.765 4.26 3.765 3.285 2.615 3.285 2.615 3.685 2.385 3.685  ;
        POLYGON 6.285 1.655 10.965 1.655 10.965 0.68 14.555 0.68 14.555 1.64 14.325 1.64 14.325 0.91 11.195 0.91 11.195 1.885 6.515 1.885 6.515 2.115 6.285 2.115  ;
        POLYGON 13.665 1.315 13.895 1.315 13.895 1.87 14.985 1.87 14.985 1.315 15.215 1.315 15.215 1.87 16.155 1.87 16.155 3.215 15.925 3.215 15.925 2.1 14.315 2.1 14.315 3.215 14.085 3.215 14.085 2.115 13.665 2.115  ;
        POLYGON 12.545 1.315 13.295 1.315 13.295 3.455 18.46 3.455 18.46 2.415 18.69 2.415 18.69 3.685 13.065 3.685 13.065 1.655 12.545 1.655  ;
        POLYGON 17.965 2.885 18 2.885 18 1.97 16.735 1.97 16.735 2.115 16.505 2.115 16.505 1.74 18.905 1.74 18.905 1.315 19.135 1.315 19.135 1.975 19.475 1.975 19.475 2.315 18.91 2.315 18.91 2.025 18.23 2.025 18.23 3.225 17.965 3.225  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1
