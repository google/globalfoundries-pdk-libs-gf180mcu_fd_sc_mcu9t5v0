# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__tieh
  CLASS core gf180mcu_fd_sc_mcu9t5v0__tiehIGH ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__tieh 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 2.24 BY 5.04 ;
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 2.89 1.53 2.89 1.53 3.7 1.27 3.7  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.25 4.59 0.25 2.945 0.48 2.945 0.48 4.59 1.6 4.59 2.24 4.59 2.24 5.49 1.6 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 2.24 -0.45 2.24 0.45 0.48 0.45 0.48 1.355 0.25 1.355 0.25 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.875 1.83 1.37 1.83 1.37 1.315 1.6 1.315 1.6 2.06 0.875 2.06  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__tieh
