# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__and4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.16 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.115 2.165 0.975 2.165 0.975 2.71 0.115 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.23 1.21 2.09 1.21 2.09 2.115 1.23 2.115  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.32 1.21 3.21 1.21 3.21 2.115 2.32 2.115  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.716 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.83 2.33 4.5 2.33 4.5 2.71 3.83 2.71  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.19 2.89 5.235 2.89 5.585 2.89 5.585 0.845 6.045 0.845 6.045 3.685 5.235 3.685 5.19 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.305 4.59 0.305 3.155 0.535 3.155 0.535 4.59 2.345 4.59 2.345 3.155 2.575 3.155 2.575 4.59 4.565 4.59 4.565 4.345 4.795 4.345 4.795 4.59 5.235 4.59 6.16 4.59 6.16 5.49 5.235 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 6.16 -0.45 6.16 0.45 4.795 0.45 4.795 1.35 4.565 1.35 4.565 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.325 2.695 3.595 2.695 3.595 2.985 4.73 2.985 4.73 2.005 3.44 2.005 3.44 0.98 0.535 0.98 0.535 1.355 0.305 1.355 0.305 0.75 3.67 0.75 3.67 1.775 5.235 1.775 5.235 2.115 4.96 2.115 4.96 3.215 3.365 3.215 3.365 2.925 1.555 2.925 1.555 3.215 1.325 3.215  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_1
