# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nor4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.77 4.33 1.77 4.33 2.555 4.07 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 2.27 3.26 2.27 3.26 2.71 2.92 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 2.27 2.14 2.27 2.14 2.71 1.8 2.71  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.311 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.71 0.71 2.71  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.4916 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.68 1.595 0.68 1.595 1.21 3.605 1.21 3.605 0.68 3.835 0.68 3.835 2.785 4.855 2.785 4.855 4.36 4.625 4.36 4.625 3.015 3.51 3.015 3.51 1.44 1.365 1.44  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 5.6 4.59 5.6 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 4.955 0.45 4.955 1.005 4.725 1.005 4.725 0.45 2.715 0.45 2.715 0.98 2.485 0.98 2.485 0.45 0.475 0.45 0.475 1.005 0.245 1.005 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor4_1
