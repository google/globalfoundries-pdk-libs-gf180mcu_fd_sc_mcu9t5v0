# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.6 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 1.21 4.89 1.21 4.89 2.115 4.63 2.115  ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.235 1.505 2.235 1.505 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.125 2.875 16.885 2.875 17.115 2.875 17.115 1.655 15.285 1.655 15.285 0.845 15.515 0.845 15.515 1.395 17.51 1.395 17.51 0.815 17.77 0.815 17.77 3.685 17.165 3.685 17.165 3.105 16.885 3.105 15.355 3.105 15.355 3.685 15.125 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.31 4.59 1.31 3.95 1.65 3.95 1.65 4.59 3.185 4.59 3.185 3.905 3.415 3.905 3.415 4.59 6.035 4.59 7.125 4.59 7.125 3.045 7.355 3.045 7.355 4.59 8.175 4.59 8.855 4.59 12.065 4.59 12.065 3.875 12.295 3.875 12.295 4.59 12.79 4.59 14.105 4.59 14.105 3.875 14.335 3.875 14.335 4.59 16.145 4.59 16.145 3.875 16.375 3.875 16.375 4.59 16.885 4.59 18.185 4.59 18.185 3.875 18.415 3.875 18.415 4.59 19.6 4.59 19.6 5.49 16.885 5.49 12.79 5.49 8.855 5.49 8.175 5.49 6.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.6 -0.45 19.6 0.45 18.875 0.45 18.875 1.165 18.645 1.165 18.645 0.45 16.635 0.45 16.635 1.165 16.405 1.165 16.405 0.45 14.395 0.45 14.395 1.165 14.165 1.165 14.165 0.45 12.155 0.45 12.155 1.165 11.925 1.165 11.925 0.45 7.52 0.45 7.52 0.625 7.29 0.625 7.29 0.45 3.435 0.45 3.435 1.435 3.205 1.435 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 3.425 1.805 3.425 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.445 6.035 3.445 6.035 4.315 5.805 4.315 5.805 3.675 0.575 3.675 0.575 4.235 0.345 4.235  ;
        POLYGON 5.165 1.315 5.395 1.315 5.395 2.415 8.175 2.415 8.175 2.755 5.395 2.755 5.395 3.215 5.165 3.215  ;
        POLYGON 6.685 1.775 8.625 1.775 8.625 1.315 8.855 1.315 8.855 3.685 8.62 3.685 8.62 2.115 6.685 2.115  ;
        POLYGON 2.385 2.525 3.845 2.525 3.845 1.895 2.485 1.895 2.485 1.315 2.715 1.315 2.715 1.665 3.845 1.665 3.845 0.69 5.89 0.69 5.89 0.855 9.01 0.855 9.01 0.69 10.855 0.69 10.855 2.755 10.625 2.755 10.625 1.085 5.665 1.085 5.665 0.92 4.075 0.92 4.075 2.755 2.615 2.755 2.615 3.215 2.385 3.215  ;
        POLYGON 9.745 1.315 9.975 1.315 9.975 3.455 11.705 3.455 11.705 2.47 12.79 2.47 12.79 2.7 11.935 2.7 11.935 3.685 9.745 3.685  ;
        POLYGON 11.265 1.775 13.045 1.775 13.045 0.845 13.31 0.845 13.31 1.975 16.885 1.975 16.885 2.315 13.315 2.315 13.315 3.685 13.085 3.685 13.085 2.115 11.265 2.115  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffq_4
