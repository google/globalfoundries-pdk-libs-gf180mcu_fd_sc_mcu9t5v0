* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__oai33_2 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(((A1 + A2) + A3) * ((B1 + B2) + B3))
M_i_5_0 VSS B3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_1 net_0 B2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_1 VSS B1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3_0 net_0 B1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_0 VSS B2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_5_1 net_0 B3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 ZN A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 ZN A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_0 A3 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_11_0 net_4_0 B3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_1 net_3_0 B2 net_4_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_1 ZN B1 net_3_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0 net_3_1 B1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_10_0 net_4_1 B2 net_3_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11_1 VDD B3 net_4_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0 net_2_0 A3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 net_1_0 A2 net_2_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_1 ZN A1 net_1_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0 net_1_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 net_2_1 A2 net_1_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_1 VDD A3 net_2_1 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
