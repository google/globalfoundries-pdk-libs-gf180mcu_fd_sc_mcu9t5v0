# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtn_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtn_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.64 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.35 1.77 11.675 1.77 11.675 2.71 11.35 2.71  ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 1.77 2.65 1.77 2.65 2.71 2.39 2.71  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.4716 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.275 0.815 16.65 0.815 16.65 4.21 16.275 4.21  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.435 4.59 1.435 3.4 1.665 3.4 1.665 4.59 2.715 4.59 5.805 4.59 5.805 3.4 6.035 3.4 6.035 4.59 8.345 4.59 8.625 4.59 8.625 3.4 8.855 3.4 8.855 4.59 9.35 4.59 12.025 4.59 12.025 3.4 12.255 3.4 12.255 4.59 12.695 4.59 15.255 4.59 15.255 3.4 15.485 3.4 15.485 4.59 15.98 4.59 17.295 4.59 17.295 3.4 17.525 3.4 17.525 4.59 17.92 4.59 17.92 5.49 15.98 5.49 12.695 5.49 9.35 5.49 8.345 5.49 2.715 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 17.675 0.45 17.675 1.625 17.445 1.625 17.445 0.45 15.435 0.45 15.435 1.625 15.205 1.625 15.205 0.45 14.395 0.45 14.395 1.155 14.165 1.155 14.165 0.45 12.155 0.45 12.155 1.155 11.925 1.155 11.925 0.45 8.755 0.45 8.755 1.155 8.525 1.155 8.525 0.45 5.795 0.45 5.795 1.155 5.565 1.155 5.565 0.45 1.65 0.45 1.65 1.1 1.31 1.1 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.815 0.475 0.815 0.475 1.31 1.16 1.31 1.16 1.33 2.065 1.33 2.065 0.815 2.715 0.815 2.715 1.155 2.295 1.155 2.295 1.56 1.065 1.56 1.065 1.54 0.245 1.54  ;
        POLYGON 3.39 1.845 6.685 1.845 6.685 0.815 7.055 0.815 7.055 3.9 6.825 3.9 6.825 2.075 4.775 2.075 4.775 2.71 4.435 2.71 4.435 2.075 3.39 2.075  ;
        POLYGON 3.16 2.835 4.24 2.835 4.24 2.94 6.495 2.94 6.495 4.13 8.115 4.13 8.115 1.885 8.345 1.885 8.345 4.36 6.265 4.36 6.265 3.17 4.275 3.17 4.275 4.21 4.045 4.21 4.045 3.065 2.93 3.065 2.93 1.385 3.605 1.385 3.605 0.815 3.835 0.815 3.835 1.615 3.16 1.615  ;
        POLYGON 7.405 0.815 7.635 0.815 7.635 1.425 8.805 1.425 8.805 1.94 9.35 1.94 9.35 2.17 8.575 2.17 8.575 1.655 7.835 1.655 7.835 3.9 7.405 3.9  ;
        POLYGON 10.535 2.91 11.235 2.91 11.235 3.72 11.005 3.72 11.005 3.14 10.305 3.14 10.305 1.31 11.09 1.31 11.09 1.54 10.535 1.54  ;
        POLYGON 9.645 0.815 9.875 0.815 9.875 3.98 11.565 3.98 11.565 2.94 12.465 2.94 12.465 2.415 12.695 2.415 12.695 3.17 11.795 3.17 11.795 4.21 9.645 4.21  ;
        POLYGON 12.99 1.31 13.33 1.31 13.33 1.33 14.015 1.33 14.015 1.94 15.98 1.94 15.98 2.17 14.015 2.17 14.015 4.21 13.785 4.21 13.785 1.56 12.99 1.56  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtn_2
