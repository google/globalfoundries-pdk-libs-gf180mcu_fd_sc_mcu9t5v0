# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 24.64 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.07 1.77 4.33 1.77 4.33 2.03 4.835 2.03 4.835 2.37 4.33 2.37 4.33 2.71 4.07 2.71  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 1.77 0.415 1.77 0.415 2.71 0.15 2.71  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.03 2.035 2.03 2.035 2.37 0.97 2.37 0.97 2.71 0.71 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.19 1.77 5.625 1.77 5.625 2.71 5.19 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.46815 ;
    PORT
      LAYER METAL1 ;
        POLYGON 20.705 0.845 20.935 0.845 20.935 1.92 22.55 1.92 22.55 1.21 22.945 1.21 22.945 0.845 23.175 0.845 23.175 1.655 22.81 1.655 22.81 2.15 20.935 2.15 20.935 3.415 23.035 3.415 23.035 4.25 22.805 4.25 22.805 3.645 20.985 3.645 20.985 4.25 20.705 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.465 4.59 10.52 4.59 11.095 4.59 13.085 4.59 13.085 3.44 13.315 3.44 13.315 4.59 14.435 4.59 17.645 4.59 17.645 3.55 17.875 3.55 17.875 4.59 18.44 4.59 19.735 4.59 19.735 3.875 19.965 3.875 19.965 4.59 20.255 4.59 21.775 4.59 21.775 3.875 22.005 3.875 22.005 4.59 23.93 4.59 23.93 3.875 24.16 3.875 24.16 4.59 24.64 4.59 24.64 5.49 20.255 5.49 18.44 5.49 14.435 5.49 11.095 5.49 10.52 5.49 3.055 5.49 0 5.49 0 4.59 1.645 4.59 1.645 3.44 1.875 3.44 1.875 4.59 3.055 4.59 5.235 4.59 5.235 3.905 8.17 3.905 8.17 4.135 5.465 4.135  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 24.64 -0.45 24.64 0.45 24.295 0.45 24.295 1.165 24.065 1.165 24.065 0.45 22.055 0.45 22.055 1.165 21.825 1.165 21.825 0.45 19.815 0.45 19.815 1.6 19.585 1.6 19.585 0.45 17.975 0.45 17.975 1.395 17.745 1.395 17.745 0.45 13.15 0.45 13.15 0.625 12.92 0.625 12.92 0.45 7.795 0.45 7.795 0.625 7.565 0.625 7.565 0.45 5.735 0.45 5.735 0.625 5.505 0.625 5.505 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.625 2.98 2.825 2.98 2.825 1.535 0.245 1.535 0.245 0.79 0.475 0.79 0.475 1.305 3.055 1.305 3.055 3.21 0.855 3.21 0.855 4.25 0.625 4.25  ;
        POLYGON 6.865 2.875 8.225 2.875 8.225 1.655 6.225 1.655 6.225 1.315 8.455 1.315 8.455 3.215 6.865 3.215  ;
        POLYGON 3.325 0.79 3.555 0.79 3.555 0.855 9.855 0.855 9.855 1.435 9.625 1.435 9.625 1.085 3.555 1.085 3.555 1.13 3.325 1.13  ;
        POLYGON 3.405 3.44 3.635 3.44 3.635 3.445 10.52 3.445 10.52 3.785 10.29 3.785 10.29 3.675 3.635 3.675 3.635 4.25 3.405 4.25  ;
        POLYGON 8.905 1.315 9.135 1.315 9.135 2.03 11.095 2.03 11.095 2.37 9.135 2.37 9.135 3.215 8.905 3.215  ;
        POLYGON 10.745 1.315 11.54 1.315 11.54 1.57 13.755 1.57 13.755 2.37 13.525 2.37 13.525 1.8 11.555 1.8 11.555 4.25 11.325 4.25 11.325 1.655 10.745 1.655  ;
        POLYGON 12.645 2.03 12.875 2.03 12.875 2.6 14.205 2.6 14.205 1.315 14.435 1.315 14.435 4.25 14.205 4.25 14.205 2.83 12.645 2.83  ;
        POLYGON 11.37 0.69 11.71 0.69 11.71 0.855 14.73 0.855 14.73 0.69 16.125 0.69 16.125 2.86 15.785 2.86 15.785 1.085 11.37 1.085  ;
        POLYGON 15.325 1.315 15.555 1.315 15.555 3.09 17.665 3.09 17.665 2.085 18.44 2.085 18.44 2.315 17.895 2.315 17.895 3.32 15.555 3.32 15.555 4.25 15.325 4.25  ;
        POLYGON 17.205 1.625 18.865 1.625 18.865 0.79 19.095 0.79 19.095 2.03 20.255 2.03 20.255 2.37 18.965 2.37 18.965 4.25 18.735 4.25 18.735 1.855 17.435 1.855 17.435 2.37 17.205 2.37  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_4
