# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__and3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.2 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.245 1.73 3.115 1.73 3.115 2.15 1.245 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.79 2.38 3.995 2.38 3.995 1.77 5 1.77 5 2.61 1.79 2.61  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 2.33 0.995 2.33 0.995 2.84 5.785 2.84 5.785 2.415 6.02 2.415 6.02 3.07 0.15 3.07  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER METAL1 ;
        POLYGON 7.55 2.925 9.26 2.925 9.58 2.925 9.58 1.6 7.25 1.6 7.25 0.895 9.93 0.895 9.93 3.63 9.26 3.63 7.55 3.63  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.505 0.475 3.505 0.475 4.59 2.285 4.59 2.285 3.975 2.515 3.975 2.515 4.59 4.325 4.59 4.325 3.975 4.555 3.975 4.555 4.59 6.585 4.59 6.585 3.875 6.815 3.875 6.815 4.59 8.625 4.59 8.625 3.875 8.855 3.875 8.855 4.59 9.26 4.59 10.665 4.59 10.665 3.875 10.895 3.875 10.895 4.59 11.2 4.59 11.2 5.49 9.26 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 11.2 -0.45 11.2 0.45 10.895 0.45 10.895 1.165 10.665 1.165 10.665 0.45 8.71 0.45 8.71 0.64 8.37 0.64 8.37 0.45 6.415 0.45 6.415 1.165 6.185 1.165 6.185 0.45 0.555 0.45 0.555 0.695 0.325 0.695 0.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.265 3.3 6.625 3.3 6.625 1.625 5.5 1.625 5.5 1.52 3.305 1.52 3.305 0.71 3.535 0.71 3.535 1.29 5.755 1.29 5.755 1.395 6.855 1.395 6.855 1.97 9.26 1.97 9.26 2.31 6.855 2.31 6.855 3.53 5.575 3.53 5.575 4.11 5.345 4.11 5.345 3.53 3.535 3.53 3.535 4.11 3.305 4.11 3.305 3.53 1.495 3.53 1.495 4.11 1.265 4.11  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_4
