# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 13.44 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 1.77 1.02 1.77 1.02 2.06 0.41 2.06 0.41 2.71 0.15 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.13 1.83 6.07 1.83 6.07 2.65 5.13 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.2448 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.11 2.965 11.075 2.965 11.585 2.965 11.585 1.62 9.18 1.62 9.18 0.73 9.63 0.73 9.63 1.39 11.64 1.39 11.64 0.73 11.87 0.73 11.87 3.9 11.19 3.9 11.19 3.31 11.075 3.31 9.41 3.31 9.41 3.9 9.11 3.9  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 3.845 1.545 3.845 1.545 4.59 6.04 4.59 6.04 3.8 6.27 3.8 6.27 4.59 8.13 4.59 8.13 3.88 8.36 3.88 8.36 4.59 10.17 4.59 10.17 3.88 10.4 3.88 10.4 4.59 11.075 4.59 12.21 4.59 12.21 3.09 12.44 3.09 12.44 4.59 13.44 4.59 13.44 5.49 11.075 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 13.44 -0.45 13.44 0.45 12.99 0.45 12.99 1.54 12.76 1.54 12.76 0.45 10.75 0.45 10.75 1.16 10.52 1.16 10.52 0.45 8.51 0.45 8.51 0.69 8.28 0.69 8.28 0.45 6.325 0.45 6.325 0.635 5.985 0.635 5.985 0.45 1.595 0.45 1.595 1.07 1.365 1.07 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.295 3.09 1.25 3.09 1.25 1.54 0.245 1.54 0.245 0.73 0.475 0.73 0.475 1.31 1.48 1.31 1.48 1.83 2.09 1.83 2.09 2.29 3.595 2.29 3.595 2.755 3.365 2.755 3.365 2.52 1.86 2.52 1.86 2.06 1.48 2.06 1.48 3.32 0.525 3.32 0.525 3.9 0.295 3.9  ;
        POLYGON 5.02 2.88 6.53 2.88 6.53 1.595 4.865 1.595 4.865 1.365 6.76 1.365 6.76 3.11 5.25 3.11 5.25 3.9 5.02 3.9  ;
        POLYGON 2.485 0.73 3.315 0.73 3.315 0.905 7.445 0.905 7.445 1.04 8.95 1.04 8.95 1.85 10.265 1.85 10.265 2.11 8.72 2.11 8.72 1.27 7.235 1.27 7.235 1.135 3.32 1.135 3.32 1.83 4.175 1.83 4.175 3.9 3.945 3.9 3.945 2.06 3.09 2.06 3.09 0.96 2.715 0.96 2.715 1.54 2.485 1.54  ;
        POLYGON 2.925 3.09 3.155 3.09 3.155 4.13 4.405 4.13 4.405 1.6 3.55 1.6 3.55 1.37 4.635 1.37 4.635 4.13 5.58 4.13 5.58 3.34 7.115 3.34 7.115 2.505 11.075 2.505 11.075 2.735 7.345 2.735 7.345 4.15 7.11 4.15 7.11 3.57 5.81 3.57 5.81 4.36 2.925 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_4
