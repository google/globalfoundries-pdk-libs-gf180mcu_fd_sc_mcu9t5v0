# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.84 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 2.27 4.01 2.27 4.01 2.5 3.77 2.5 3.77 2.71 2.945 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.04 2.33 17.275 2.33 17.275 2.71 16.04 2.71  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.22 1.77 15.115 1.77 15.115 2.15 14.22 2.15  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 2.2 1.575 2.2 1.575 2.71 0.685 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.245 0.845 20.57 0.845 20.57 3.685 20.245 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.425 1.495 3.425 1.495 4.59 2.035 4.59 3.005 4.59 3.005 3.515 3.235 3.515 3.235 4.59 4.835 4.59 7.305 4.59 7.305 4.49 7.535 4.49 7.535 4.59 10.505 4.59 10.505 4.49 10.735 4.49 10.735 4.59 12.55 4.59 14.39 4.59 14.39 3.95 14.73 3.95 14.73 4.59 16.43 4.59 16.43 3.95 16.77 3.95 16.77 4.59 18.195 4.59 18.525 4.59 18.525 3.425 18.755 3.425 18.755 4.59 19.245 4.59 19.245 3.875 19.475 3.875 19.475 4.59 19.795 4.59 21.285 4.59 21.285 3.875 21.515 3.875 21.515 4.59 21.84 4.59 21.84 5.49 19.795 5.49 18.195 5.49 12.55 5.49 4.835 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.84 -0.45 21.84 0.45 21.595 0.45 21.595 1.165 21.365 1.165 21.365 0.45 19.355 0.45 19.355 1.165 19.125 1.165 19.125 0.45 16.635 0.45 16.635 1.225 16.405 1.225 16.405 0.45 8.875 0.45 8.875 1.425 8.645 1.425 8.645 0.45 3.515 0.45 3.515 1.425 3.285 1.425 3.285 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.94 1.805 2.94 1.805 1.74 0.245 1.74 0.245 1.315 0.475 1.315 0.475 1.51 2.035 1.51 2.035 3.17 0.475 3.17 0.475 3.75 0.245 3.75  ;
        POLYGON 4.025 2.73 4.405 2.73 4.405 1.315 4.635 1.315 4.635 2.96 4.255 2.96 4.255 3.685 4.025 3.685  ;
        POLYGON 2.285 1.315 2.715 1.315 2.715 3.055 3.695 3.055 3.695 3.975 4.835 3.975 4.835 4.315 3.465 4.315 3.465 3.285 2.515 3.285 2.515 3.685 2.285 3.685  ;
        POLYGON 6.065 3.35 8.775 3.35 8.775 3.8 6.065 3.8  ;
        POLYGON 5.045 2.875 5.525 2.875 5.525 1.315 5.755 1.315 5.755 2.875 9.325 2.875 9.325 2.575 9.555 2.575 9.555 3.105 5.275 3.105 5.275 3.685 5.045 3.685  ;
        POLYGON 9.265 3.46 10.605 3.46 10.605 2.345 7.035 2.345 7.035 2.455 6.805 2.455 6.805 2.115 10.605 2.115 10.605 1.315 10.835 1.315 10.835 3.57 11.685 3.57 11.685 2.875 11.915 2.875 11.915 3.8 9.265 3.8  ;
        POLYGON 5.57 4.03 12.55 4.03 12.55 4.26 5.57 4.26  ;
        POLYGON 5.985 1.655 10.145 1.655 10.145 0.68 13.79 0.68 13.79 0.91 10.375 0.91 10.375 1.885 6.215 1.885 6.215 2.115 5.985 2.115  ;
        POLYGON 12.845 1.2 15.68 1.2 15.68 2.875 15.695 2.875 15.695 3.215 15.45 3.215 15.45 1.54 13.955 1.54 13.955 3.215 13.725 3.215 13.725 1.65 12.845 1.65  ;
        POLYGON 11.725 1.315 11.955 1.315 11.955 1.88 12.935 1.88 12.935 3.455 17.965 3.455 17.965 2.415 18.195 2.415 18.195 3.685 12.705 3.685 12.705 2.11 11.725 2.11  ;
        POLYGON 15.91 1.87 18.365 1.87 18.365 1.315 18.595 1.315 18.595 1.775 19.795 1.775 19.795 2.115 17.735 2.115 17.735 3.215 17.505 3.215 17.505 2.1 15.91 2.1  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2
