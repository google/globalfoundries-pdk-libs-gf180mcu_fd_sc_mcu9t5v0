# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__addf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 23.52 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.7 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.705 1.86 6.785 1.86 6.785 2.71 5.705 2.71  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.7 ;
    PORT
      LAYER METAL1 ;
        POLYGON 16.965 2.33 18.53 2.33 18.53 2.71 16.965 2.71  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.525 ;
    PORT
      LAYER METAL1 ;
        POLYGON 7.33 1.92 8.11 1.92 11.415 1.92 11.91 1.92 11.91 1.77 12.17 1.77 12.17 1.92 15.495 1.92 15.99 1.92 15.99 2.15 15.495 2.15 11.415 2.15 8.11 2.15 7.33 2.15  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER METAL1 ;
        POLYGON 19.635 2.875 20.725 2.875 20.725 1.655 19.685 1.655 19.685 0.845 19.915 0.845 19.915 1.425 21.925 1.425 21.925 0.845 22.155 0.845 22.155 1.655 21.185 1.655 21.185 2.875 22.105 2.875 22.105 3.685 21.875 3.685 21.875 3.105 19.865 3.105 19.865 3.685 19.635 3.685  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.81585 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.84 2.875 4.015 2.875 4.015 3.685 3.785 3.685 3.785 3.105 1.675 3.105 1.675 3.685 1.445 3.685 1.445 2.875 2.38 2.875 2.38 1.655 1.445 1.655 1.445 0.845 1.675 0.845 1.675 1.425 3.685 1.425 3.685 0.845 3.915 0.845 3.915 1.655 2.84 1.655  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.325 4.59 0.325 3.875 0.555 3.875 0.555 4.59 2.555 4.59 2.555 3.875 2.785 3.875 2.785 4.59 4.905 4.59 4.905 3.875 5.135 3.875 5.135 4.59 8.11 4.59 10.065 4.59 10.065 3.905 10.295 3.905 10.295 4.59 11.37 4.59 12.205 4.59 12.205 3.435 12.435 3.435 12.435 4.59 14.145 4.59 14.145 3.435 14.375 3.435 14.375 4.59 15.395 4.59 18.465 4.59 18.465 3.875 18.695 3.875 18.695 4.59 19.235 4.59 20.75 4.59 20.75 3.875 20.98 3.875 20.98 4.59 22.945 4.59 22.945 3.875 23.175 3.875 23.175 4.59 23.52 4.59 23.52 5.49 19.235 5.49 15.395 5.49 11.37 5.49 8.11 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 23.52 -0.45 23.52 0.45 23.275 0.45 23.275 1.165 23.045 1.165 23.045 0.45 21.035 0.45 21.035 1.165 20.805 1.165 20.805 0.45 18.795 0.45 18.795 1.165 18.565 1.165 18.565 0.45 14.375 0.45 14.375 1.215 14.145 1.215 14.145 0.45 12.535 0.45 12.535 1.215 12.305 1.215 12.305 0.45 10.295 0.45 10.295 1.215 10.065 1.215 10.065 0.45 5.035 0.45 5.035 1.165 4.805 1.165 4.805 0.45 2.795 0.45 2.795 1.165 2.565 1.165 2.565 0.45 0.555 0.45 0.555 1.165 0.325 1.165 0.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 4.31 1.83 5.245 1.83 5.245 1.315 8.11 1.315 8.11 1.545 5.475 1.545 5.475 2.94 7.825 2.94 7.825 2.875 8.055 2.875 8.055 3.685 7.825 3.685 7.825 3.17 5.245 3.17 5.245 2.06 4.595 2.06 4.595 2.585 4.31 2.585  ;
        POLYGON 9.045 2.93 11.37 2.93 11.37 3.16 9.275 3.16 9.275 3.74 9.045 3.74  ;
        POLYGON 8.945 1.315 9.175 1.315 9.175 1.445 11.185 1.445 11.185 1.315 11.415 1.315 11.415 1.675 8.945 1.675  ;
        POLYGON 13.125 2.93 15.395 2.93 15.395 3.74 15.165 3.74 15.165 3.16 13.355 3.16 13.355 3.74 13.125 3.74  ;
        POLYGON 13.025 1.315 13.255 1.315 13.255 1.445 15.265 1.445 15.265 1.315 15.495 1.315 15.495 1.675 13.025 1.675  ;
        POLYGON 8.45 2.47 15.855 2.47 15.855 2.94 19.005 2.94 19.005 2.005 16.385 2.005 16.385 1.315 16.615 1.315 16.615 1.775 19.235 1.775 19.235 3.17 16.515 3.17 16.515 3.75 16.285 3.75 16.285 3.17 15.625 3.17 15.625 2.7 8.45 2.7  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_4
