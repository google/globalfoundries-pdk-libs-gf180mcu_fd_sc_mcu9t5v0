# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai221_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.32 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.53 2.215 7.76 2.215 7.76 2.89 9.075 2.89 9.075 2.27 11.14 2.27 11.14 2.5 9.305 2.5 9.305 3.27 7.53 3.27  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.99 1.77 8.25 1.77 8.25 2.215 8.845 2.215 8.845 2.555 7.99 2.555  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 2.15 3.21 2.15 3.21 2.71 2.95 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 1.83 2.165 1.83 2.165 2.325 2.5 2.325 2.5 2.94 4.575 2.94 4.575 2.215 5.425 2.215 5.425 2.555 4.805 2.555 4.805 3.17 2.27 3.17 2.27 2.555 1.21 2.555  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 3.35 2.125 3.35 2.125 3.4 5.035 3.4 5.035 2.785 6.16 2.785 6.395 2.785 6.395 2.215 6.625 2.215 6.625 3.015 6.16 3.015 5.265 3.015 5.265 3.63 1.98 3.63 1.98 3.58 0.71 3.58  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.2165 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.295 3.81 1.835 3.81 1.835 3.86 5.495 3.86 5.495 3.55 6.16 3.55 10.79 3.55 10.79 2.89 11.435 2.89 11.435 1.985 8.48 1.985 8.48 1.54 8.12 1.54 8.12 1.31 8.71 1.31 8.71 1.755 10.415 1.755 10.415 1.14 10.645 1.14 10.645 1.755 11.665 1.755 11.665 3.78 7.205 3.78 7.205 4.36 6.975 4.36 6.975 3.78 6.16 3.78 5.725 3.78 5.725 4.09 3.765 4.09 3.765 4.36 3.535 4.36 3.535 4.09 1.69 4.09 1.69 4.04 0.525 4.04 0.525 4.36 0.295 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 4.27 1.545 4.27 1.545 4.59 5.955 4.59 5.955 4.02 6.16 4.02 6.185 4.02 6.185 4.59 9.245 4.59 9.245 4.02 9.475 4.02 9.475 4.59 11.765 4.59 12.32 4.59 12.32 5.49 11.765 5.49 6.16 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.32 -0.45 12.32 0.45 5.04 0.45 5.04 0.64 4.7 0.64 4.7 0.45 2.8 0.45 2.8 0.64 2.46 0.64 2.46 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.34 1.33 6.16 1.33 6.16 1.56 1.34 1.56  ;
        POLYGON 0.245 0.715 0.475 0.715 0.475 0.87 7.055 0.87 7.055 0.68 11.765 0.68 11.765 1.525 11.535 1.525 11.535 0.91 9.525 0.91 9.525 1.525 9.295 1.525 9.295 0.91 7.285 0.91 7.285 1.19 7.055 1.19 7.055 1.1 0.475 1.1 0.475 1.525 0.245 1.525  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai221_2
