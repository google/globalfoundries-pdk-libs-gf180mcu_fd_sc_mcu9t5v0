# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.72 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.885 2.065 2.115 2.065 2.115 2.58 3.28 2.58 3.51 2.58 3.51 2.12 4.4 2.12 4.4 2.35 3.77 2.35 3.77 2.81 3.28 2.81 1.885 2.81  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.81 2.12 1.435 2.12 1.435 3.04 3.28 3.04 4.43 3.04 4.43 2.89 4.66 2.89 4.66 2.12 5.47 2.12 5.47 2.35 4.89 2.35 4.89 3.27 3.28 3.27 1.205 3.27 1.205 2.35 0.81 2.35  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.675 3.5 5.305 3.5 5.305 2.58 5.75 2.58 5.75 1.37 4.69 1.37 4.69 1.14 6.01 1.14 6.01 2.81 5.535 2.81 5.535 3.73 3.905 3.73 3.905 4.31 3.675 4.31  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.285 4.59 0.285 3.5 0.515 3.5 0.515 4.59 2.325 4.59 2.325 3.5 2.555 3.5 2.555 4.59 3.28 4.59 5.765 4.59 5.765 3.5 5.995 3.5 5.995 4.59 6.15 4.59 6.72 4.59 6.72 5.49 6.15 5.49 3.28 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 6.72 -0.45 6.72 0.45 2.555 0.45 2.555 1.355 2.325 1.355 2.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.285 1.015 0.515 1.015 0.515 1.605 2.575 1.605 2.575 2.12 3.28 2.12 3.28 2.35 2.345 2.35 2.345 1.835 0.515 1.835 0.515 2.58 0.975 2.58 0.975 3.5 1.535 3.5 1.535 4.31 1.305 4.31 1.305 3.73 0.745 3.73 0.745 2.81 0.285 2.81  ;
        POLYGON 3.625 0.68 6.15 0.68 6.15 0.91 3.855 0.91 3.855 1.655 3.625 1.655  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor2_1
