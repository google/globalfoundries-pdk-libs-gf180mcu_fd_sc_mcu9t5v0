# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 13.44 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.335 1.77 3.335 2.71 2.95 2.71  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 2.275 1.37 2.275 1.37 1.31 4.175 1.31 4.175 1.77 5.495 1.77 5.495 2.56 5.265 2.56 5.265 2.15 4.175 2.15 4.175 2.56 3.945 2.56 3.945 1.54 1.6 1.54 1.6 2.505 0.705 2.505  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.34 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.495 1.77 2.495 2.71 1.83 2.71  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.55 1.77 8.875 1.77 8.875 2.71 8.55 2.71  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.425 0.845 12.735 0.845 12.735 4.21 12.425 4.21  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.4 1.495 3.4 1.495 4.59 3.065 4.59 3.065 3.89 3.295 3.89 3.295 4.59 6.645 4.59 6.645 3.89 6.875 3.89 6.875 4.59 7.315 4.59 8.925 4.59 8.925 3.4 9.155 3.4 9.155 4.59 11.225 4.59 11.225 3.43 11.455 3.43 11.455 4.59 11.915 4.59 13.44 4.59 13.44 5.49 11.915 5.49 7.315 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 13.44 -0.45 13.44 0.45 11.615 0.45 11.615 1.165 11.385 1.165 11.385 0.45 7.47 0.45 7.47 1.075 7.13 1.075 7.13 0.45 1.595 0.45 1.595 1.08 1.365 1.08 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.79 0.475 0.79 0.475 2.94 4.545 2.94 4.545 2.38 4.775 2.38 4.775 3.17 0.475 3.17 0.475 4.21 0.245 4.21  ;
        POLYGON 2.045 3.4 7.085 3.4 7.085 3.02 5.725 3.02 5.725 1.13 4.385 1.13 4.385 0.79 5.955 0.79 5.955 2.79 7.315 2.79 7.315 3.63 5.055 3.63 5.055 4.21 4.825 4.21 4.825 3.63 2.275 3.63 2.275 4.21 2.045 4.21  ;
        POLYGON 7.905 2.94 9.325 2.94 9.325 1.54 6.415 1.54 6.415 2.56 6.185 2.56 6.185 1.31 9.325 1.31 9.325 0.79 9.555 0.79 9.555 2.22 10.715 2.22 10.715 2.56 9.555 2.56 9.555 3.17 8.135 3.17 8.135 4.21 7.905 4.21  ;
        POLYGON 10.205 2.97 11.685 2.97 11.685 1.655 10.045 1.655 10.045 1.315 10.275 1.315 10.275 1.425 11.915 1.425 11.915 3.2 10.435 3.2 10.435 4.21 10.205 4.21  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_1
