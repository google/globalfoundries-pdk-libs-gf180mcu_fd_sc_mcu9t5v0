# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.88 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.19 1.77 5.645 1.77 5.645 2.71 5.19 2.71  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.9952 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.465 2.965 11.365 2.965 12.03 2.965 12.265 2.965 12.265 1.6 10.025 1.6 10.025 0.79 10.255 0.79 10.255 1.37 12.265 1.37 12.265 0.84 12.495 0.84 12.495 3.195 12.03 3.195 11.735 3.195 11.735 4.21 11.505 4.21 11.505 3.195 11.365 3.195 9.93 3.195 9.93 4.21 9.465 4.21  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.37 4.59 1.37 3.845 1.6 3.845 1.6 4.59 6.045 4.59 6.045 4.28 6.275 4.28 6.275 4.59 8.265 4.59 8.265 3.4 8.495 3.4 8.495 4.59 10.485 4.59 10.485 3.88 10.715 3.88 10.715 4.59 11.365 4.59 12.03 4.59 12.88 4.59 12.88 5.49 12.03 5.49 11.365 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 12.88 -0.45 12.88 0.45 11.375 0.45 11.375 1.02 11.145 1.02 11.145 0.45 8.955 0.45 8.955 1.16 8.725 1.16 8.725 0.45 6.575 0.45 6.575 0.62 6.235 0.62 6.235 0.45 1.65 0.45 1.65 1.02 1.42 1.02 1.42 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.35 2.94 3.335 2.94 3.335 2.06 1.2 2.06 1.2 1.54 0.3 1.54 0.3 0.68 0.53 0.68 0.53 1.31 1.43 1.31 1.43 1.83 3.565 1.83 3.565 3.17 0.58 3.17 0.58 4.21 0.35 4.21  ;
        POLYGON 5.025 2.94 6.75 2.94 6.75 1.54 4.92 1.54 4.92 1.31 7.09 1.31 7.09 2.06 6.98 2.06 6.98 3.17 5.255 3.17 5.255 3.75 5.025 3.75  ;
        POLYGON 2.895 3.4 3.125 3.4 3.125 3.98 4.375 3.98 4.375 1.655 4.255 1.655 4.255 1.315 4.605 1.315 4.605 3.98 5.605 3.98 5.605 3.82 7.245 3.82 7.245 2.505 11.365 2.505 11.365 2.735 7.475 2.735 7.475 4.05 5.825 4.05 5.825 4.21 2.895 4.21  ;
        POLYGON 2.54 0.68 2.77 0.68 2.77 0.85 7.835 0.85 7.835 1.83 12.03 1.83 12.03 2.06 7.605 2.06 7.605 1.08 4.025 1.08 4.025 2.94 4.145 2.94 4.145 3.75 3.795 3.75 3.795 1.49 2.54 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_3
