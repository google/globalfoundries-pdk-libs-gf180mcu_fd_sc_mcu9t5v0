* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I B:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(((A1 + A2) * B) * C)
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_0 net_1_0 B net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_0 VSS C net_1_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_1 net_1_1 C VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_1 net_0 B net_1_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_5_1 net_2_0 A2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_4_1 ZN A1 net_2_0 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_4_0 net_2_1 A1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_5_0 VDD A2 net_2_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_0 ZN B VDD VNW pfet_05v0 W=1.460000U L=0.500000U
M_i_7_0 VDD C ZN VNW pfet_05v0 W=1.460000U L=0.500000U
M_i_7_1 ZN C VDD VNW pfet_05v0 W=1.460000U L=0.500000U
M_i_6_1 VDD B ZN VNW pfet_05v0 W=1.460000U L=0.500000U
.ENDS
