# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyc_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyc_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.14 0.99 1.14 0.99 1.84 0.65 1.84  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.565 2.875 11.995 2.875 12.225 2.875 12.225 1.655 10.565 1.655 10.565 0.845 10.795 0.845 10.795 1.425 12.47 1.425 12.47 0.845 13.035 0.845 13.035 1.655 12.455 1.655 12.455 2.875 12.935 2.875 12.935 3.685 12.705 3.685 12.705 3.105 11.995 3.105 10.795 3.105 10.795 3.685 10.565 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.71 1.495 3.71 1.495 4.59 4.315 4.59 4.665 4.59 4.665 3.71 4.895 3.71 4.895 4.59 8.315 4.59 8.665 4.59 8.665 3.71 8.895 3.71 8.895 4.59 11.585 4.59 11.585 3.875 11.815 3.875 11.815 4.59 11.995 4.59 13.825 4.59 13.825 3.875 14.055 3.875 14.055 4.59 14.56 4.59 14.56 5.49 11.995 5.49 8.315 5.49 4.315 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 14.155 0.45 14.155 1.165 13.925 1.165 13.925 0.45 11.915 0.45 11.915 1.165 11.685 1.165 11.685 0.45 8.995 0.45 8.995 0.935 8.765 0.935 8.765 0.45 4.995 0.45 4.995 0.935 4.765 0.935 4.765 0.45 1.595 0.45 1.595 0.965 1.365 0.965 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.53 1.87 2.53 1.87 2.06 2.21 2.06 2.21 2.76 0.475 2.76 0.475 4.05 0.19 4.05 0.19 0.68 0.53 0.68 0.53 0.91 0.42 0.91  ;
        POLYGON 1.485 2.99 4.085 2.99 4.085 1.715 1.43 1.715 1.43 1.485 4.315 1.485 4.315 3.33 1.485 3.33  ;
        POLYGON 4.665 1.315 4.995 1.315 4.995 1.83 6.21 1.83 6.21 2.53 5.87 2.53 5.87 2.06 4.895 2.06 4.895 3.33 4.665 3.33  ;
        POLYGON 5.485 2.76 8.085 2.76 8.085 1.6 5.43 1.6 5.43 1.37 8.315 1.37 8.315 2.99 5.715 2.99 5.715 3.33 5.485 3.33  ;
        POLYGON 8.665 1.315 8.995 1.315 8.995 1.975 11.995 1.975 11.995 2.315 8.895 2.315 8.895 3.33 8.665 3.33  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyc_4
