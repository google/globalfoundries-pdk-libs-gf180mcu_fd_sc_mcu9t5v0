# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__and3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.16 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.115 2.15 0.97 2.15 0.97 2.71 0.115 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.21 2.15 2.09 2.15 2.09 2.71 1.21 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.39 2.29 3.21 2.29 3.21 2.71 2.39 2.71  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.48 0.845 4.89 0.845 4.89 3.685 4.48 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.32 4.59 1.32 3.875 1.55 3.875 1.55 4.59 3.36 4.59 3.36 3.875 3.59 3.875 3.59 4.59 4.21 4.59 5.58 4.59 5.58 3.875 5.81 3.875 5.81 4.59 6.16 4.59 6.16 5.49 4.21 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 6.16 -0.45 6.16 0.45 5.83 0.45 5.83 1.165 5.6 1.165 5.6 0.45 3.59 0.45 3.59 1.165 3.36 1.165 3.36 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 3.3 3.98 3.3 3.98 1.92 0.3 1.92 0.3 0.845 0.53 0.845 0.53 1.69 4.21 1.69 4.21 3.53 2.57 3.53 2.57 4.11 2.34 4.11 2.34 3.53 0.245 3.53  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_2
