* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__fillcap_16 VDD VNW VPW VSS
*.PININFO VDD:P VNW:P VPW:P VSS:G
M_i_17 net_3 net_2 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23 net_4 net_5 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_24 net_7 net_9 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_17_23_55 net_6 net_8 VSS VPW nmos_5p0 W=1.320000U L=1.000000U
M_i_19 VDD net_3 net_2 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7 VDD net_4 net_5 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_33 VDD net_7 net_9 VNW pmos_5p0 W=1.830000U L=1.000000U
M_i_19_7_23 VDD net_6 net_8 VNW pmos_5p0 W=1.830000U L=1.000000U
.ENDS
