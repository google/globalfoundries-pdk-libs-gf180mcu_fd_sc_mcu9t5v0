# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__or4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.27 1.07 2.27 1.07 2.71 0.71 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.555 1.83 2.555  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.39 2.27 3.26 2.27 3.26 2.71 2.39 2.71  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.51 2.27 4.38 2.27 4.38 2.71 3.51 2.71  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7295 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.75 2.89 6.025 2.89 6.025 0.68 6.255 0.68 6.255 4.36 5.75 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 4.675 4.59 4.675 3.55 4.905 3.55 4.905 4.59 5.625 4.59 7.045 4.59 7.045 3.55 7.275 3.55 7.275 4.59 7.84 4.59 7.84 5.49 5.625 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 7.375 0.45 7.375 1.49 7.145 1.49 7.145 0.45 4.955 0.45 4.955 1.02 4.725 1.02 4.725 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.02 0.245 1.02 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 3.09 4.61 3.09 4.61 1.48 1.365 1.48 1.365 0.68 1.595 0.68 1.595 1.25 3.605 1.25 3.605 0.68 3.835 0.68 3.835 1.25 4.84 1.25 4.84 2.215 5.625 2.215 5.625 2.555 4.84 2.555 4.84 3.32 0.575 3.32 0.575 4.36 0.345 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_2
