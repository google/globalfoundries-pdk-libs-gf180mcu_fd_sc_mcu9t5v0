# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.33 2.09 2.33 2.09 2.71 0.87 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.735 1.77 6.115 1.77 6.115 2.15 5.735 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.2448 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.785 2.97 8.56 2.97 8.96 2.97 8.96 1.62 7.685 1.62 7.685 0.68 7.915 0.68 7.915 1.39 9.925 1.39 9.925 0.68 10.155 0.68 10.155 1.62 9.42 1.62 9.42 2.97 10.055 2.97 10.055 3.78 9.825 3.78 9.825 3.2 8.56 3.2 8.015 3.2 8.015 3.78 7.785 3.78  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.845 1.595 3.845 1.595 4.59 4.725 4.59 4.725 4.35 4.955 4.35 4.955 4.59 6.765 4.59 6.765 3.88 6.995 3.88 6.995 4.59 8.56 4.59 8.805 4.59 8.805 3.88 9.035 3.88 9.035 4.59 10.845 4.59 10.845 3.88 11.075 3.88 11.075 4.59 11.76 4.59 11.76 5.49 8.56 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 11.275 0.45 11.275 1.16 11.045 1.16 11.045 0.45 9.035 0.45 9.035 1.16 8.805 1.16 8.805 0.45 6.85 0.45 6.85 0.635 6.51 0.635 6.51 0.45 4.61 0.45 4.61 0.635 4.27 0.635 4.27 0.45 1.595 0.45 1.595 1.165 1.365 1.165 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 1.83 2.55 1.83 2.55 2.47 3.65 2.47 3.65 2.7 2.32 2.7 2.32 2.06 0.575 2.06 0.575 3.685 0.245 3.685  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.91 6.575 0.91 6.575 1.85 8.56 1.85 8.56 2.08 6.345 2.08 6.345 1.14 3.32 1.14 3.32 1.83 4.165 1.83 4.165 3.215 3.935 3.215 3.935 2.06 3.09 2.06 3.09 1.49 2.485 1.49  ;
        POLYGON 2.915 2.93 3.145 2.93 3.145 3.51 4.395 3.51 4.395 1.6 3.55 1.6 3.55 1.37 4.625 1.37 4.625 2.505 8.56 2.505 8.56 2.735 5.975 2.735 5.975 3.72 5.745 3.72 5.745 2.735 4.625 2.735 4.625 3.74 2.915 3.74  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_4
