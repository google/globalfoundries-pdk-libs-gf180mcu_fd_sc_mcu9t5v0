# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai22_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.04 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.73 1.755 13.745 1.755 13.745 2.27 15.53 2.27 15.53 2.5 13.515 2.5 13.515 1.985 11.34 1.985 11.34 2.5 10.73 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.885 2.215 10.115 2.215 10.115 2.73 12.47 2.73 12.47 2.215 13.285 2.215 13.285 2.73 17.485 2.73 17.485 2.215 17.715 2.215 17.715 2.96 9.885 2.96  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.11 1.77 5.04 1.77 5.04 2.27 6.57 2.27 6.57 2.5 4.81 2.5 4.81 2.15 4.58 2.15 4.58 2.04 3.45 2.04 3.45 2.5 3.11 2.5  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.875 2.215 1.105 2.215 1.105 2.73 4.04 2.73 4.04 2.27 4.38 2.27 4.38 2.73 6.8 2.73 6.8 2.27 8.81 2.27 8.81 2.5 7.03 2.5 7.03 2.96 0.875 2.96  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.5585 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.585 3.19 17.945 3.19 17.945 1.475 10.27 1.475 10.27 1.14 10.61 1.14 10.61 1.245 12.51 1.245 12.51 1.14 15.09 1.14 15.09 1.245 16.99 1.245 16.99 1.14 18.175 1.14 18.175 3.45 18.33 3.45 18.33 3.83 16.205 3.83 16.205 4.36 15.975 4.36 15.975 3.42 11.625 3.42 11.625 4.36 11.395 4.36 11.395 3.42 7.095 3.42 7.095 4.36 6.865 4.36 6.865 3.42 2.815 3.42 2.815 4.36 2.585 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 4.675 4.59 4.675 3.65 4.905 3.65 4.905 4.59 9.105 4.59 9.105 3.65 9.335 3.65 9.335 4.59 13.635 4.59 13.635 3.65 13.865 3.65 13.865 4.59 18.065 4.59 18.065 4.06 18.295 4.06 18.295 4.59 18.635 4.59 19.04 4.59 19.04 5.49 18.635 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 19.04 -0.45 19.04 0.45 8.315 0.45 8.315 1.07 8.085 1.07 8.085 0.45 6.075 0.45 6.075 1.07 5.845 1.07 5.845 0.45 3.835 0.45 3.835 1.07 3.605 1.07 3.605 0.45 1.595 0.45 1.595 1.07 1.365 1.07 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.73 0.475 0.73 0.475 1.31 2.485 1.31 2.485 0.73 2.715 0.73 2.715 1.31 4.725 1.31 4.725 0.73 4.955 0.73 4.955 1.31 6.965 1.31 6.965 0.73 7.195 0.73 7.195 1.31 9.205 1.31 9.205 0.68 18.635 0.68 18.635 1.54 18.405 1.54 18.405 0.91 16.21 0.91 16.21 1.015 15.87 1.015 15.87 0.91 11.73 0.91 11.73 1.015 11.39 1.015 11.39 0.91 9.435 0.91 9.435 1.54 0.245 1.54  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai22_4
