# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.412 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.65 2.215 4.205 2.215 4.205 2.65 0.65 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.2024 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.025 3.09 8.92 3.09 9.15 3.09 9.15 1.745 6.025 1.745 6.025 0.945 6.255 0.945 6.255 1.515 8.265 1.515 8.265 0.945 8.495 0.945 8.495 1.515 10.505 1.515 10.505 0.945 10.735 0.945 10.735 1.515 12.745 1.515 12.745 0.945 12.975 0.945 12.975 1.745 9.65 1.745 9.65 3.09 12.875 3.09 12.875 4.36 12.645 4.36 12.645 3.32 10.635 3.32 10.635 4.36 10.23 4.36 10.23 3.32 8.92 3.32 8.395 3.32 8.395 4.36 8.165 4.36 8.165 3.32 6.255 3.32 6.255 4.36 6.025 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.875 4.855 3.875 4.855 4.59 7.045 4.59 7.045 3.55 7.275 3.55 7.275 4.59 8.92 4.59 9.285 4.59 9.285 3.55 9.515 3.55 9.515 4.59 11.525 4.59 11.525 3.55 11.755 3.55 11.755 4.59 13.51 4.59 13.765 4.59 13.765 3.55 13.995 3.55 13.995 4.59 14.56 4.59 14.56 5.49 13.51 5.49 8.92 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 14.095 0.45 14.095 1.285 13.865 1.285 13.865 0.45 11.855 0.45 11.855 1.215 11.625 1.215 11.625 0.45 9.615 0.45 9.615 1.215 9.385 1.215 9.385 0.45 7.375 0.45 7.375 1.285 7.145 1.285 7.145 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.365 3.09 4.435 3.09 4.435 1.745 1.365 1.745 1.365 0.945 1.595 0.945 1.595 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 4.665 1.515 4.665 2.27 8.92 2.27 8.92 2.65 4.665 2.65 4.665 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
        POLYGON 9.88 2.27 13.51 2.27 13.51 2.65 9.88 2.65  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_8
