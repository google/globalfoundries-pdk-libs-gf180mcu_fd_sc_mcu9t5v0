# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.656 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.265 4.26 2.265 4.26 2.645 0.63 2.645  ;
        POLYGON 5.36 2.215 8.88 2.215 8.88 2.65 5.36 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.284 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 4.63 3.09 4.63 1.985 1.365 1.985 1.365 0.68 1.595 0.68 1.595 1.755 3.575 1.755 3.575 0.68 3.835 0.68 3.835 1.755 5.845 1.755 5.845 0.68 6.075 0.68 6.075 1.755 8.085 1.755 8.085 0.68 8.315 0.68 8.315 1.985 5.13 1.985 5.13 3.09 8.215 3.09 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 10.08 4.59 10.08 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.165 4.725 1.165 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_8
