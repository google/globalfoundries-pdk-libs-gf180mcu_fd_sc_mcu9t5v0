* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
*.PININFO A1:I A2:I A3:I Z:O VDD:P VNW:P VPW:P VSS:G
*.EQN Z=((A1 + A2) + A3)
M_i_2 VSS A1 Z_neg VPW nfet_05v0 W=0.525000U L=0.600000U
M_i_3 Z_neg A2 VSS VPW nfet_05v0 W=0.525000U L=0.600000U
M_i_4 VSS A3 Z_neg VPW nfet_05v0 W=0.525000U L=0.600000U
M_i_0 Z Z_neg VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_5 net_0 A1 Z_neg VNW pfet_05v0 W=0.915000U L=0.500000U
M_i_6 net_1 A2 net_0 VNW pfet_05v0 W=0.915000U L=0.500000U
M_i_7 VDD A3 net_1 VNW pfet_05v0 W=0.915000U L=0.500000U
M_i_1 Z Z_neg VDD VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
