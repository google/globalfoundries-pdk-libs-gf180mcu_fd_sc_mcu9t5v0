* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__inv_8 I ZN VDD VNW VPW VSS
*.PININFO I:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!I
M_i_0_0_x8_0 ZN I VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0_x8_1 VSS I ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0_x8_2 ZN I VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0_x8_3 VSS I ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0_x8_4 ZN I VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0_x8_5 VSS I ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0_x8_6 ZN I VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0_x8_7 VSS I ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_0_x8_0 ZN I VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_0_x8_1 VDD I ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_0_x8_2 ZN I VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_0_x8_3 VDD I ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_0_x8_4 ZN I VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_0_x8_5 VDD I ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_0_x8_6 ZN I VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_0_x8_7 VDD I ZN VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
