* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__latrnq_4 D E RN Q VDD VNW VPW VSS
*.PININFO D:I E:I RN:I Q:O VDD:P VNW:P VPW:P VSS:G
M_tn3 net7 E VSS VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn10 net1 RN VSS VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn9 net2 D net1 VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn8 net2 E net3 VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn7 net3 net7 net4 VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn5 net5 net0 net4 VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn0 VSS RN net5 VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn6 net0 net3 VSS VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn6_109 net0 net3 VSS VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn4 net6 net0 VSS VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn4_77 net6 net0 VSS VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn1 Q net6 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_tn1_38 Q net6 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_tn1_15 Q net6 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_tn1_38_14 Q net6 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_tp2 net7 E VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp8 VDD RN net3 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp6 net8 D VDD VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp5 net3 net7 net8 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp4 net9 E net3 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp3 net9 net0 VDD VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp9 net0 net3 VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp9_110 net0 net3 VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp7 net6 net0 VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp7_78 net6 net0 VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp0 Q net6 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_tp0_27 Q net6 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_tp0_24 Q net6 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_tp0_27_20 Q net6 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
