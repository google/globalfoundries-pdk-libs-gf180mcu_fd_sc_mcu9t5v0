# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.118 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.275 1.77 6.01 1.77 6.01 2.215 6.675 2.215 6.675 2.555 1.275 2.555  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.3036 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.485 3.09 13.205 3.09 13.465 3.09 13.465 1.54 8.485 1.54 8.485 1.18 8.715 1.18 8.715 1.31 10.725 1.31 10.725 0.74 10.955 0.74 10.955 1.31 12.965 1.31 12.965 0.74 13.195 0.74 13.195 1.31 15.205 1.31 15.205 0.74 15.435 0.74 15.435 1.31 17.445 1.31 17.445 0.74 17.675 0.74 17.675 1.31 19.685 1.31 19.685 1.18 19.915 1.18 19.915 1.54 14.35 1.54 14.35 3.09 19.815 3.09 19.815 4.36 19.585 4.36 19.585 3.32 17.575 3.32 17.575 4.36 17.345 4.36 17.345 3.32 15.335 3.32 15.335 4.36 14.71 4.36 14.71 3.32 13.205 3.32 13.095 3.32 13.095 4.36 12.865 4.36 12.865 3.32 10.855 3.32 10.855 4.36 10.625 4.36 10.625 3.32 8.715 3.32 8.715 4.36 8.485 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.465 4.59 0.465 3.55 0.695 3.55 0.695 4.59 2.605 4.59 2.605 3.55 2.835 3.55 2.835 4.59 4.845 4.59 4.845 3.55 5.075 3.55 5.075 4.59 7.365 4.59 7.365 3.875 7.595 3.875 7.595 4.59 9.505 4.59 9.505 3.55 9.735 3.55 9.735 4.59 11.745 4.59 11.745 3.55 11.975 3.55 11.975 4.59 13.205 4.59 13.985 4.59 13.985 3.55 14.215 3.55 14.215 4.59 16.225 4.59 16.225 3.55 16.455 3.55 16.455 4.59 18.465 4.59 18.465 3.55 18.695 3.55 18.695 4.59 19.98 4.59 20.705 4.59 20.705 3.55 20.935 3.55 20.935 4.59 21.28 4.59 21.28 5.49 19.98 5.49 13.205 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 21.035 0.45 21.035 1.08 20.805 1.08 20.805 0.45 18.795 0.45 18.795 1.08 18.565 1.08 18.565 0.45 16.555 0.45 16.555 1.08 16.325 1.08 16.325 0.45 14.315 0.45 14.315 1.08 14.085 1.08 14.085 0.45 12.075 0.45 12.075 1.08 11.845 1.08 11.845 0.45 9.835 0.45 9.835 1.08 9.605 1.08 9.605 0.45 7.415 0.45 7.415 1.08 7.185 1.08 7.185 0.45 5.175 0.45 5.175 1.08 4.945 1.08 4.945 0.45 2.935 0.45 2.935 1.08 2.705 1.08 2.705 0.45 0.475 0.45 0.475 1.315 0.245 1.315 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.585 3.09 6.905 3.09 6.905 1.54 1.585 1.54 1.585 1.11 1.815 1.11 1.815 1.31 3.825 1.31 3.825 1.11 4.055 1.11 4.055 1.31 6.065 1.31 6.065 1.11 6.295 1.11 6.295 1.31 7.135 1.31 7.135 2.215 13.205 2.215 13.205 2.555 7.135 2.555 7.135 3.32 6.195 3.32 6.195 4.36 5.965 4.36 5.965 3.32 3.955 3.32 3.955 4.36 3.725 4.36 3.725 3.32 1.815 3.32 1.815 4.36 1.585 4.36  ;
        POLYGON 14.58 2.215 19.98 2.215 19.98 2.555 14.58 2.555  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_12
