# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.68 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.245 1.21 2.65 1.21 2.65 2.15 2.245 2.15  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.945 1.92 2.015 1.92 2.015 2.38 2.88 2.38 2.88 1.92 3.22 1.92 3.22 2.33 3.77 2.33 3.77 2.945 4.195 2.945 4.195 3.27 3.51 3.27 3.51 2.61 1.785 2.61 1.785 2.15 0.945 2.15  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.87 1.77 7.23 1.77 7.23 2.71 6.87 2.71  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.51 3.09 11.76 3.09 11.76 0.84 11.99 0.84 11.99 1.21 14 1.21 14 0.84 14.23 0.84 14.23 1.65 13.85 1.65 13.85 2.15 13.59 2.15 13.59 1.44 11.99 1.44 11.99 3.09 13.78 3.09 13.78 4.25 13.55 4.25 13.55 3.32 11.74 3.32 11.74 4.25 11.51 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.61 4.59 1.61 3.705 1.84 3.705 1.84 4.59 3.28 4.59 5.39 4.59 5.39 3.55 5.62 3.55 5.62 4.59 7.61 4.59 7.61 3.875 7.84 3.875 7.84 4.59 8.45 4.59 8.45 3.875 8.68 3.875 8.68 4.59 9.07 4.59 10.49 4.59 10.49 3.875 10.72 3.875 10.72 4.59 11.3 4.59 12.53 4.59 12.53 3.55 12.76 3.55 12.76 4.59 14.57 4.59 14.57 3.875 14.8 3.875 14.8 4.59 15.68 4.59 15.68 5.49 11.3 5.49 9.07 5.49 3.28 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 15.68 -0.45 15.68 0.45 15.35 0.45 15.35 1.16 15.12 1.16 15.12 0.45 13.11 0.45 13.11 0.69 12.88 0.69 12.88 0.45 10.87 0.45 10.87 1.16 10.64 1.16 10.64 0.45 8.63 0.45 8.63 1.16 8.4 1.16 8.4 0.45 5.77 0.45 5.77 1.31 5.54 1.31 5.54 0.45 1.67 0.45 1.67 1.305 1.44 1.305 1.44 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.32 0.88 0.55 0.88 0.55 2.66 0.815 2.66 0.815 2.84 3.28 2.84 3.28 3.18 0.82 3.18 0.82 4.36 0.59 4.36 0.59 2.89 0.32 2.89  ;
        POLYGON 3.63 3.55 3.86 3.55 3.86 4.13 4.425 4.13 4.425 1.77 3.58 1.77 3.58 0.97 3.81 0.97 3.81 1.54 6.23 1.54 6.23 2.31 6 2.31 6 1.77 4.655 1.77 4.655 4.36 3.63 4.36  ;
        POLYGON 5.1 2 5.33 2 5.33 2.905 6.715 2.905 6.715 2.94 8.84 2.94 8.84 1.65 7.68 1.65 7.68 0.84 7.91 0.84 7.91 1.42 9.07 1.42 9.07 3.17 6.82 3.17 6.82 4.25 6.59 4.25 6.59 3.135 5.1 3.135  ;
        POLYGON 9.47 0.84 9.75 0.84 9.75 1.94 11.3 1.94 11.3 2.28 9.7 2.28 9.7 4.25 9.47 4.25  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_4
