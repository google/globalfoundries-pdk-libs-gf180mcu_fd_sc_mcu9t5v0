# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.12 BY 5.04 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.22 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.23 1.77 10.49 1.77 10.49 2.71 10.23 2.71  ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.77 2.255 1.77 2.255 2.71 1.83 2.71  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 1.21 0.41 1.21 0.41 2.27 1.19 2.27 1.19 2.5 0.15 2.5  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.2452 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.15 0.695 14.61 0.695 14.61 3.685 14.15 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.21 4.59 13.915 4.59 15.12 4.59 15.12 5.49 13.915 5.49 2.935 5.49 0 5.49 0 4.59 0.845 4.59 0.845 3.435 1.075 3.435 1.075 4.59 2.935 4.59 6.025 4.59 6.025 3.91 6.255 3.91 6.255 4.59 8.98 4.59 8.98 3.895 11.2 3.895 11.2 4.005 13.01 4.005 13.01 3.425 13.24 3.425 13.24 4.235 9.21 4.235  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 15.12 -0.45 15.12 0.45 13.49 0.45 13.49 1.015 13.26 1.015 13.26 0.45 9.49 0.45 9.49 1.035 9.26 1.035 9.26 0.45 6.015 0.45 6.015 1.13 5.785 1.13 5.785 0.45 1.87 0.45 1.87 1.075 1.53 1.075 1.53 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.19 0.75 0.87 0.75 0.87 1.305 2.705 1.305 2.705 0.79 2.935 0.79 2.935 1.535 0.64 1.535 0.64 0.98 0.19 0.98  ;
        POLYGON 3.665 1.79 3.895 1.79 3.895 2.485 4.99 2.485 4.99 2.715 3.665 2.715  ;
        POLYGON 3.435 2.945 5.22 2.945 5.22 1.755 6.37 1.755 6.37 2.27 6.75 2.27 6.75 2.5 6.14 2.5 6.14 1.985 5.45 1.985 5.45 3.175 3.595 3.175 3.595 4.245 3.205 4.245 3.205 0.845 4.11 0.845 4.11 1.075 3.435 1.075  ;
        POLYGON 7.565 2.375 8.14 2.375 8.14 0.695 8.475 0.695 8.475 3.18 8.135 3.18 8.135 2.605 7.565 2.605  ;
        POLYGON 8.715 2.27 9.77 2.27 9.77 0.75 10.665 0.75 10.665 0.98 10 0.98 10 2.95 10.515 2.95 10.515 3.18 9.77 3.18 9.77 2.5 8.715 2.5  ;
        POLYGON 5.68 2.215 5.91 2.215 5.91 3.41 6.98 3.41 6.98 1.13 6.905 1.13 6.905 0.79 7.21 0.79 7.21 3.41 10.745 3.41 10.745 2.27 12.555 2.27 12.555 2.5 10.975 2.5 10.975 3.64 7.275 3.64 7.275 4.245 7.045 4.245 7.045 3.64 5.68 3.64  ;
        POLYGON 11.99 2.875 12.785 2.875 12.785 1.035 11.1 1.035 11.1 0.695 13.015 0.695 13.015 2.27 13.915 2.27 13.915 2.5 13.015 2.5 13.015 3.105 12.22 3.105 12.22 3.685 11.99 3.685  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_1
