# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 22.4 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.39 1.77 3.99 1.77 3.99 1.21 4.33 1.21 4.33 2.15 3.39 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER METAL1 ;
        POLYGON 16.755 2.32 17.77 2.32 17.77 2.71 16.755 2.71  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER METAL1 ;
        POLYGON 15.27 1.21 15.61 1.21 15.61 2.06 15.27 2.06  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.77 1.58 1.77 1.58 2.15 0.71 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER METAL1 ;
        POLYGON 20.67 0.845 21.13 0.845 21.13 3.83 20.67 3.83  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.47 4.59 1.47 3.425 1.7 3.425 1.7 4.59 2.14 4.59 3.21 4.59 3.21 3.595 3.44 3.595 3.44 4.59 7.69 4.59 7.69 4.48 7.92 4.48 7.92 4.59 10.83 4.59 10.83 4.48 11.06 4.48 11.06 4.59 12.795 4.59 14.775 4.59 14.775 3.96 15.115 3.96 15.115 4.59 16.815 4.59 16.815 3.96 17.155 3.96 17.155 4.59 18.69 4.59 18.91 4.59 18.91 3.905 19.14 3.905 19.14 4.59 19.65 4.59 19.65 3.875 19.88 3.875 19.88 4.59 20.32 4.59 21.69 4.59 21.69 3.875 21.92 3.875 21.92 4.59 22.4 4.59 22.4 5.49 20.32 5.49 18.69 5.49 12.795 5.49 2.14 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 22.4 -0.45 22.4 0.45 22.02 0.45 22.02 1.165 21.79 1.165 21.79 0.45 19.78 0.45 19.78 1.165 19.55 1.165 19.55 0.45 17.1 0.45 17.1 1.225 16.87 1.225 16.87 0.45 9.215 0.45 9.215 1.37 8.875 1.37 8.875 0.45 3.67 0.45 3.67 1.425 3.44 1.425 3.44 0.45 1.755 0.45 1.755 1.045 1.415 1.045 1.415 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.45 2.875 1.91 2.875 1.91 1.54 0.35 1.54 0.35 1.19 0.58 1.19 0.58 1.31 2.14 1.31 2.14 3.105 0.68 3.105 0.68 3.685 0.45 3.685  ;
        POLYGON 4.23 2.955 4.56 2.955 4.56 1.315 4.79 1.315 4.79 3.185 4.46 3.185 4.46 3.765 4.23 3.765  ;
        POLYGON 6.52 2.98 6.75 2.98 6.75 3.45 9.16 3.45 9.16 3.79 6.52 3.79  ;
        POLYGON 5.25 2.52 5.68 2.52 5.68 1.315 5.91 1.315 5.91 2.52 10.09 2.52 10.09 2.505 10.32 2.505 10.32 2.845 10.09 2.845 10.09 2.75 5.48 2.75 5.48 3.765 5.25 3.765  ;
        POLYGON 9.65 2.98 9.88 2.98 9.88 3.075 10.55 3.075 10.55 2.275 10.005 2.275 10.005 2.29 7.1 2.29 7.1 1.95 7.33 1.95 7.33 2.06 9.92 2.06 9.92 2.045 11.21 2.045 11.21 1.315 11.44 1.315 11.44 2.225 12.3 2.225 12.3 3.775 12.07 3.775 12.07 2.455 10.78 2.455 10.78 3.305 9.88 3.305 9.88 3.79 9.65 3.79  ;
        POLYGON 2.49 1.19 2.82 1.19 2.82 2.985 3.9 2.985 3.9 4.02 12.795 4.02 12.795 4.35 12.455 4.35 12.455 4.25 5.975 4.25 5.975 4.34 3.67 4.34 3.67 3.215 2.49 3.215  ;
        POLYGON 6.36 1.49 7.73 1.49 7.73 1.6 9.605 1.6 9.605 0.68 14.38 0.68 14.38 0.91 9.835 0.91 9.835 1.83 7.53 1.83 7.53 1.72 6.59 1.72 6.59 2.115 6.36 2.115  ;
        POLYGON 13.45 1.14 14.81 1.14 14.81 0.75 16.08 0.75 16.08 3.225 15.85 3.225 15.85 0.98 15.04 0.98 15.04 1.37 14.34 1.37 14.34 3.305 14.11 3.305 14.11 1.48 13.45 1.48  ;
        POLYGON 12.33 1.315 12.56 1.315 12.56 1.67 13.32 1.67 13.32 3.545 14.495 3.545 14.495 3.5 18.46 3.5 18.46 2.425 18.69 2.425 18.69 3.73 14.635 3.73 14.635 3.775 13.09 3.775 13.09 1.9 12.33 1.9  ;
        POLYGON 17.89 2.91 18 2.91 18 2.09 16.375 2.09 16.375 1.86 18.83 1.86 18.83 1.315 19.06 1.315 19.06 1.775 20.32 1.775 20.32 2.115 18.23 2.115 18.23 3.25 17.89 3.25  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2
