# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__addf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 16.8 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.396 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.265 2.33 3.455 2.33 3.455 2.71 2.265 2.71  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.396 ;
    PORT
      LAYER METAL1 ;
        POLYGON 13.525 2.265 13.85 2.265 13.85 2.71 13.525 2.71  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.547 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.89 2.115 7.975 2.115 11.91 2.115 11.91 1.77 12.11 1.77 12.17 1.77 12.17 2.115 12.55 2.115 12.55 2.345 12.11 2.345 7.975 2.345 3.89 2.345  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 15.83 2.89 16.145 2.89 16.145 0.845 16.475 0.845 16.475 3.685 15.83 3.685  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.3244 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 0.845 0.575 0.845 0.575 3.83 0.15 3.83  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.875 1.595 3.875 1.595 4.59 4.615 4.59 6.625 4.59 6.625 3.61 6.855 3.61 6.855 4.59 7.93 4.59 8.665 4.59 8.665 3.14 8.895 3.14 8.895 4.59 10.705 4.59 10.705 3.505 10.935 3.505 10.935 4.59 11.955 4.59 15.125 4.59 15.125 3.875 15.355 3.875 15.355 4.59 15.795 4.59 16.8 4.59 16.8 5.49 15.795 5.49 11.955 5.49 7.93 5.49 4.615 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 16.8 -0.45 16.8 0.45 15.355 0.45 15.355 1.165 15.125 1.165 15.125 0.45 10.935 0.45 10.935 1.425 10.705 1.425 10.705 0.45 9.095 0.45 9.095 1.425 8.865 1.425 8.865 0.45 6.855 0.45 6.855 1.425 6.625 1.425 6.625 0.45 1.595 0.45 1.595 1.305 1.365 1.305 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 2.035 2.94 4.615 2.94 4.615 3.79 4.385 3.79 4.385 3.17 1.805 3.17 1.805 2.06 0.87 2.06 0.87 1.655 4.385 1.655 4.385 1.315 4.615 1.315 4.615 1.885 2.035 1.885  ;
        POLYGON 5.605 3.035 7.93 3.035 7.93 3.265 5.835 3.265 5.835 3.845 5.605 3.845  ;
        POLYGON 5.505 1.315 5.735 1.315 5.735 1.655 7.745 1.655 7.745 1.315 7.975 1.315 7.975 1.885 5.505 1.885  ;
        POLYGON 9.685 3.035 11.955 3.035 11.955 3.845 11.725 3.845 11.725 3.265 9.915 3.265 9.915 3.845 9.685 3.845  ;
        POLYGON 9.585 1.315 9.815 1.315 9.815 1.655 11.45 1.655 11.45 1.31 12.11 1.31 12.11 1.54 11.68 1.54 11.68 1.885 9.585 1.885  ;
        POLYGON 5.01 2.575 13.075 2.575 13.075 2.94 14.08 2.94 14.08 2.005 12.945 2.005 12.945 1.315 13.175 1.315 13.175 1.775 15.795 1.775 15.795 2.115 14.31 2.115 14.31 3.17 13.075 3.17 13.075 3.685 12.845 3.685 12.845 2.805 5.01 2.805  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_1
