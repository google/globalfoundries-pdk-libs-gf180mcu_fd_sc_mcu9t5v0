# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.97 4.59 1.765 4.59 1.765 3.55 1.995 3.55 1.995 4.59 3.21 4.59 4.005 4.59 4.005 3.55 4.235 3.55 4.235 4.59 5.45 4.59 6.245 4.59 6.245 3.55 6.475 3.55 6.475 4.59 7.69 4.59 8.485 4.59 8.485 3.55 8.715 3.55 8.715 4.59 9.93 4.59 10.725 4.59 10.725 3.55 10.955 3.55 10.955 4.59 12.17 4.59 12.965 4.59 12.965 3.55 13.195 3.55 13.195 4.59 14.41 4.59 15.205 4.59 15.205 3.55 15.435 3.55 15.435 4.59 16.65 4.59 17.445 4.59 17.445 3.55 17.675 3.55 17.675 4.59 17.92 4.59 17.92 5.49 17.675 5.49 16.65 5.49 15.435 5.49 14.41 5.49 13.195 5.49 12.17 5.49 10.955 5.49 9.93 5.49 8.715 5.49 7.69 5.49 6.475 5.49 5.45 5.49 4.235 5.49 3.21 5.49 1.995 5.49 0.97 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 16.155 0.45 16.155 1.49 15.925 1.49 15.925 0.45 13.915 0.45 13.915 1.49 13.685 1.49 13.685 0.45 11.675 0.45 11.675 1.49 11.445 1.49 11.445 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 1.83 0.97 1.83 0.97 2.06 0.475 2.06 0.475 4.36 0.245 4.36  ;
        POLYGON 1.325 1.26 1.765 1.26 1.765 0.68 1.995 0.68 1.995 1.49 1.555 1.49 1.555 2.755 1.325 2.755  ;
        POLYGON 2.485 1.83 3.21 1.83 3.21 2.06 2.715 2.06 2.715 4.36 2.485 4.36  ;
        POLYGON 3.565 1.26 4.005 1.26 4.005 0.68 4.235 0.68 4.235 1.49 3.795 1.49 3.795 2.755 3.565 2.755  ;
        POLYGON 4.725 1.83 5.45 1.83 5.45 2.06 4.955 2.06 4.955 4.36 4.725 4.36  ;
        POLYGON 5.805 1.26 6.245 1.26 6.245 0.68 6.475 0.68 6.475 1.49 6.035 1.49 6.035 2.755 5.805 2.755  ;
        POLYGON 6.965 1.83 7.69 1.83 7.69 2.06 7.195 2.06 7.195 4.36 6.965 4.36  ;
        POLYGON 8.045 1.26 8.485 1.26 8.485 0.68 8.715 0.68 8.715 1.49 8.275 1.49 8.275 2.755 8.045 2.755  ;
        POLYGON 9.205 1.83 9.93 1.83 9.93 2.06 9.435 2.06 9.435 4.36 9.205 4.36  ;
        POLYGON 10.285 1.26 10.725 1.26 10.725 0.68 10.955 0.68 10.955 1.49 10.515 1.49 10.515 2.755 10.285 2.755  ;
        POLYGON 11.445 1.83 12.17 1.83 12.17 2.06 11.675 2.06 11.675 4.36 11.445 4.36  ;
        POLYGON 12.525 1.26 12.965 1.26 12.965 0.68 13.195 0.68 13.195 1.49 12.755 1.49 12.755 2.755 12.525 2.755  ;
        POLYGON 13.685 1.83 14.41 1.83 14.41 2.06 13.915 2.06 13.915 4.36 13.685 4.36  ;
        POLYGON 14.765 1.26 15.205 1.26 15.205 0.68 15.435 0.68 15.435 1.49 14.995 1.49 14.995 2.755 14.765 2.755  ;
        POLYGON 15.925 1.83 16.65 1.83 16.65 2.06 16.155 2.06 16.155 4.36 15.925 4.36  ;
        POLYGON 17.005 1.26 17.445 1.26 17.445 0.68 17.675 0.68 17.675 1.49 17.235 1.49 17.235 2.755 17.005 2.755  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_32
