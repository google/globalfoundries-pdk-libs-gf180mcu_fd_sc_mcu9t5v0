# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.16 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 4.03 1.77 4.03 2.15 2.95 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.97 1.83 14.655 1.83 14.655 2.17 12.97 2.17  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.33 1.53 2.33 1.53 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.19 0.845 19.45 0.845 19.45 3.685 19.19 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.305 4.59 3.305 3.145 3.535 3.145 3.535 4.59 5.15 4.59 7.525 4.59 7.525 3.96 7.755 3.96 7.755 4.59 10.005 4.59 10.005 4.005 10.235 4.005 10.235 4.59 11.575 4.59 13.985 4.59 13.985 3.145 14.215 3.145 14.215 4.59 15.235 4.59 16.025 4.59 16.025 3.615 16.255 3.615 16.255 4.59 18.185 4.59 18.185 3.875 18.415 3.875 18.415 4.59 18.855 4.59 20.16 4.59 20.16 5.49 18.855 5.49 15.235 5.49 11.575 5.49 5.15 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 20.16 -0.45 20.16 0.45 18.315 0.45 18.315 1.165 18.085 1.165 18.085 0.45 16.475 0.45 16.475 1.265 16.245 1.265 16.245 0.45 7.635 0.45 7.635 1.245 7.405 1.245 7.405 0.45 3.435 0.45 3.435 1.245 3.205 1.245 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.325 1.135 4.555 1.135 4.555 3.785 4.325 3.785  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 2.685 3.995 2.685 3.995 4.13 5.15 4.13 5.15 4.36 3.765 4.36 3.765 2.915 2.615 2.915 2.615 3.685 2.385 3.685  ;
        POLYGON 5.445 1.135 5.675 1.135 5.675 2.11 8.47 2.11 8.47 2.34 5.675 2.34 5.675 3.785 5.445 3.785  ;
        POLYGON 6.07 1.65 7.865 1.65 7.865 0.68 10.51 0.68 10.51 0.91 8.095 0.91 8.095 1.88 6.07 1.88  ;
        POLYGON 6.81 2.57 9.785 2.57 9.785 1.315 10.015 1.315 10.015 2.975 11.135 2.975 11.135 3.315 8.765 3.315 8.765 2.8 6.81 2.8  ;
        POLYGON 5.97 3.5 8.035 3.5 8.035 3.545 11.575 3.545 11.575 4.315 11.345 4.315 11.345 3.775 7.895 3.775 7.895 3.73 6.31 3.73 6.31 4.36 5.97 4.36  ;
        POLYGON 12.74 2.4 13.495 2.4 13.495 2.685 15.235 2.685 15.235 3.785 15.005 3.785 15.005 2.915 13.495 2.915 13.495 3.685 13.265 3.685 13.265 2.63 12.51 2.63 12.51 1.655 12.025 1.655 12.025 1.26 14.215 1.26 14.215 1.6 12.74 1.6  ;
        POLYGON 10.905 0.8 15.115 0.8 15.115 1.83 16.97 1.83 16.97 2.06 14.885 2.06 14.885 1.03 11.135 1.03 11.135 1.885 12.155 1.885 12.155 3.685 11.925 3.685 11.925 2.115 10.905 2.115  ;
        POLYGON 15.585 2.515 17.365 2.515 17.365 1.315 17.595 1.315 17.595 2.39 18.855 2.39 18.855 2.73 17.455 2.73 17.455 3.215 15.585 3.215  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_1
