* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 I Z VDD VNW VPW VSS
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nmos_5p0 W=0.550000U L=0.600000U
M_i_2_1 VSS I Z_neg VPW nmos_5p0 W=0.550000U L=0.600000U
M_i_0_0 Z Z_neg VSS VPW nmos_5p0 W=0.600000U L=0.600000U
M_i_0_1 VSS Z_neg Z VPW nmos_5p0 W=0.600000U L=0.600000U
M_i_0_2 Z Z_neg VSS VPW nmos_5p0 W=0.600000U L=0.600000U
M_i_0_3 VSS Z_neg Z VPW nmos_5p0 W=0.600000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pmos_5p0 W=1.375000U L=0.500000U
M_i_3_1 VDD I Z_neg VNW pmos_5p0 W=1.375000U L=0.500000U
M_i_1_0 Z Z_neg VDD VNW pmos_5p0 W=1.375000U L=0.500000U
M_i_1_1 VDD Z_neg Z VNW pmos_5p0 W=1.375000U L=0.500000U
M_i_1_2 Z Z_neg VDD VNW pmos_5p0 W=1.375000U L=0.500000U
M_i_1_3 VDD Z_neg Z VNW pmos_5p0 W=1.375000U L=0.500000U
.ENDS
