# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 31.92 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.545 2.33 1.575 2.33 1.575 2.71 0.545 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.536 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.3 2.15 12.125 2.15 12.125 2.71 5.3 2.71  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 12.9792 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.52 3.365 27.62 3.365 27.775 3.365 28.53 3.365 28.53 1.635 14.595 1.635 14.595 0.865 30.505 0.865 30.505 1.65 29.09 1.65 29.09 4.175 27.775 4.175 27.62 4.175 14.52 4.175  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.505 4.59 1.505 3.845 1.735 3.845 1.735 4.59 4.86 4.59 4.86 4.37 5.2 4.37 5.2 4.59 6.9 4.59 6.9 4.37 7.24 4.37 7.24 4.59 8.94 4.59 8.94 4.37 9.28 4.37 9.28 4.59 11.28 4.59 11.28 4.37 11.62 4.37 11.62 4.59 13.5 4.59 13.5 4.405 13.84 4.405 13.84 4.59 15.54 4.59 15.54 4.405 15.88 4.405 15.88 4.59 17.58 4.59 17.58 4.405 17.92 4.405 17.92 4.59 19.62 4.59 19.62 4.405 19.96 4.405 19.96 4.59 21.66 4.59 21.66 4.405 22 4.405 22 4.59 23.7 4.59 23.7 4.405 24.04 4.405 24.04 4.59 25.74 4.59 25.74 4.405 26.08 4.405 26.08 4.59 27.62 4.59 27.775 4.59 27.78 4.59 27.78 4.405 28.12 4.405 28.12 4.59 29.875 4.59 29.875 3.88 30.105 3.88 30.105 4.59 31.92 4.59 31.92 5.49 27.775 5.49 27.62 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 31.92 -0.45 31.92 0.45 31.625 0.45 31.625 1.16 31.395 1.16 31.395 0.45 29.44 0.45 29.44 0.635 29.1 0.635 29.1 0.45 27.2 0.45 27.2 0.635 26.86 0.635 26.86 0.45 24.96 0.45 24.96 0.635 24.62 0.635 24.62 0.45 22.72 0.45 22.72 0.635 22.38 0.635 22.38 0.45 20.48 0.45 20.48 0.635 20.14 0.635 20.14 0.45 18.24 0.45 18.24 0.635 17.9 0.635 17.9 0.45 16 0.45 16 0.635 15.66 0.635 15.66 0.45 13.78 0.45 13.78 0.635 13.405 0.635 13.405 0.45 11.52 0.45 11.52 0.635 11.18 0.635 11.18 0.45 9.28 0.45 9.28 0.635 8.94 0.635 8.94 0.45 7.04 0.45 7.04 0.635 6.7 0.635 6.7 0.45 4.61 0.45 4.61 0.625 4.27 0.625 4.27 0.45 1.595 0.45 1.595 0.695 1.365 0.695 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.485 2.94 1.805 2.94 1.805 1.6 0.19 1.6 0.19 1.37 2.035 1.37 2.035 2.94 3.365 2.94 3.365 2.415 3.595 2.415 3.595 3.17 0.715 3.17 0.715 3.75 0.485 3.75  ;
        POLYGON 2.925 3.445 4.405 3.445 4.405 1.655 3.605 1.655 3.605 1.315 4.635 1.315 4.635 3.33 12.355 3.33 12.355 2.47 27.62 2.47 27.62 2.755 12.7 2.755 12.7 4.14 2.925 4.14  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.855 5.865 0.855 5.865 0.865 14.145 0.865 14.145 1.865 27.775 1.865 27.775 2.16 13.855 2.16 13.855 1.65 5.635 1.65 5.635 1.085 3.375 1.085 3.375 1.955 4.175 1.955 4.175 3.215 3.945 3.215 3.945 2.185 3.145 2.185 3.145 1.49 2.485 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_16
