# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__addh_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.03 2.27 3.84 2.27 3.84 2.94 5.75 2.94 5.75 2.27 7.16 2.27 7.16 2.5 6.01 2.5 6.01 3.17 3.61 3.17 3.61 2.5 3.03 2.5  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.07 2.15 4.33 2.15 4.33 2.71 4.07 2.71  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.27 0.77 1.615 0.77 1.615 4.355 1.27 4.355  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7295 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.985 0.77 10.49 0.77 10.49 1.59 10.215 1.59 10.215 4.355 9.985 4.355  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.315 4.59 0.315 3.875 0.545 3.875 0.545 4.59 2.455 4.59 2.455 3.875 2.685 3.875 2.685 4.59 4.545 4.59 4.545 3.875 4.775 3.875 4.775 4.59 5.365 4.59 5.365 3.875 5.595 3.875 5.595 4.59 8.865 4.59 8.865 3.875 9.095 3.875 9.095 4.59 9.635 4.59 11.055 4.59 11.055 3.875 11.285 3.875 11.285 4.59 11.76 4.59 11.76 5.49 9.635 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 11.335 0.45 11.335 1.58 11.105 1.58 11.105 0.45 9.095 0.45 9.095 1.58 8.865 1.58 8.865 0.45 2.735 0.45 2.735 1.58 2.505 1.58 2.505 0.45 0.495 0.45 0.495 1.58 0.265 1.58 0.265 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 5.265 0.68 7.735 0.68 7.735 1.11 7.505 1.11 7.505 0.91 5.495 0.91 5.495 1.58 5.265 1.58  ;
        POLYGON 2.015 1.855 2.245 1.855 2.245 2.385 2.8 2.385 2.8 3.4 7.945 3.4 7.945 2.04 4.545 2.04 4.545 0.77 4.775 0.77 4.775 1.81 8.175 1.81 8.175 3.63 3.755 3.63 3.755 4.325 3.525 4.325 3.525 3.63 2.57 3.63 2.57 2.665 2.015 2.665  ;
        POLYGON 7.505 3.875 8.405 3.875 8.405 1.57 6.385 1.57 6.385 1.14 6.615 1.14 6.615 1.34 8.635 1.34 8.635 2.27 9.4 2.27 9.4 1.835 9.635 1.835 9.635 2.645 8.635 2.645 8.635 4.215 7.505 4.215  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_2
