# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 25.76 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.21 1.77 3.21 2.2 4.075 2.2 4.075 2.43 3.21 2.43 3.21 2.71 2.95 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.898 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.43 1.77 21.795 1.77 21.795 2.71 21.43 2.71  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.41 1.77 0.41 2.145 0.94 2.145 0.94 2.71 0.15 2.71  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.745 1.77 20.01 1.77 20.01 2.71 19.745 2.71  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.71 1.83 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 2.33 7.13 2.33 7.13 2.71 6.31 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 24.775 2.33 25.285 2.33 25.285 0.845 25.515 0.845 25.515 2.56 25.05 2.56 25.05 4.075 24.775 4.075  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.34 4.59 1.34 3.435 1.57 3.435 1.57 4.59 5.11 4.59 5.11 3.905 5.34 3.905 5.34 4.59 7.03 4.59 7.03 4.005 7.37 4.005 7.37 4.59 9.075 4.59 9.515 4.59 12.125 4.59 12.125 4.33 12.355 4.33 12.355 4.59 15.245 4.59 15.245 4.505 15.475 4.505 15.475 4.59 17.21 4.59 19.275 4.59 19.275 4.07 19.505 4.07 19.505 4.59 21.48 4.59 21.48 4.265 21.82 4.265 21.82 4.59 23.245 4.59 23.575 4.59 23.575 3.74 23.805 3.74 23.805 4.59 24.425 4.59 25.76 4.59 25.76 5.49 24.425 5.49 23.245 5.49 17.21 5.49 9.515 5.49 9.075 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 25.76 -0.45 25.76 0.45 24.395 0.45 24.395 1.6 24.165 1.6 24.165 0.45 21.31 0.45 21.31 1.08 20.97 1.08 20.97 0.45 13.655 0.45 13.655 1.425 13.425 1.425 13.425 0.45 7.615 0.45 7.615 1.135 7.385 1.135 7.385 0.45 5.76 0.45 5.76 0.535 5.53 0.535 5.53 0.45 1.675 0.45 1.675 1.08 1.335 1.08 1.335 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.32 2.94 2.49 2.94 2.49 1.54 0.27 1.54 0.27 0.795 0.5 0.795 0.5 1.31 2.72 1.31 2.72 2.94 4.73 2.94 4.73 2.145 4.96 2.145 4.96 3.17 0.55 3.17 0.55 4.075 0.32 4.075  ;
        POLYGON 6.065 2.94 7.525 2.94 7.525 2.055 6.265 2.055 6.265 1.225 6.495 1.225 6.495 1.825 7.755 1.825 7.755 3.28 6.065 3.28  ;
        POLYGON 3.35 3.435 5.73 3.435 5.73 3.545 8.845 3.545 8.845 2.965 9.075 2.965 9.075 3.775 5.53 3.775 5.53 3.665 3.58 3.665 3.58 4.245 3.35 4.245  ;
        POLYGON 3.35 0.765 6.955 0.765 6.955 1.365 8.045 1.365 8.045 0.765 9.455 0.765 9.455 1.425 9.225 1.425 9.225 0.995 8.275 0.995 8.275 1.595 6.725 1.595 6.725 0.995 3.58 0.995 3.58 1.135 3.35 1.135  ;
        POLYGON 8.105 2.255 8.505 2.255 8.505 1.225 8.735 1.225 8.735 2.145 9.515 2.145 9.515 2.485 8.335 2.485 8.335 3.27 8.105 3.27  ;
        POLYGON 10.885 3.265 13.555 3.265 13.555 3.605 10.885 3.605  ;
        POLYGON 9.865 2.895 10.345 2.895 10.345 1.085 10.575 1.085 10.575 2.715 14.485 2.715 14.485 2.605 14.715 2.605 14.715 2.945 10.57 2.945 10.57 3.125 10.095 3.125 10.095 3.945 9.865 3.945  ;
        POLYGON 14.045 3.265 14.945 3.265 14.945 2.375 12.095 2.375 12.095 2.485 11.865 2.485 11.865 2.145 15.905 2.145 15.905 1.315 16.715 1.315 16.715 3.895 16.485 3.895 16.485 1.545 16.135 1.545 16.135 2.375 15.175 2.375 15.175 3.605 14.045 3.605  ;
        POLYGON 10.39 3.87 15.825 3.87 15.825 4.125 17.21 4.125 17.21 4.355 15.65 4.355 15.65 4.275 15.42 4.275 15.42 4.1 10.73 4.1 10.73 4.35 10.39 4.35  ;
        POLYGON 10.925 1.655 15.445 1.655 15.445 0.68 18.835 0.68 18.835 2.485 18.605 2.485 18.605 0.91 15.675 0.91 15.675 1.885 11.155 1.885 11.155 2.485 10.925 2.485  ;
        POLYGON 18.145 1.315 18.375 1.315 18.375 2.715 19.065 2.715 19.065 0.795 19.295 0.795 19.295 1.31 20.525 1.31 20.525 3.77 20.295 3.77 20.295 1.54 19.295 1.54 19.295 2.945 18.755 2.945 18.755 3.31 18.525 3.31 18.525 2.945 18.145 2.945  ;
        POLYGON 17.025 1.315 17.735 1.315 17.735 3.61 19.965 3.61 19.965 4 20.61 4 20.61 3.985 21.025 3.985 21.025 3.76 23.015 3.76 23.015 2.145 23.245 2.145 23.245 3.99 21.255 3.99 21.255 4.215 20.695 4.215 20.695 4.23 19.735 4.23 19.735 3.84 17.735 3.84 17.735 3.95 17.505 3.95 17.505 1.655 17.025 1.655  ;
        POLYGON 20.82 1.31 23.445 1.31 23.445 0.795 23.69 0.795 23.69 1.83 24.425 1.83 24.425 2.485 24.195 2.485 24.195 2.06 23.46 2.06 23.46 1.54 22.785 1.54 22.785 3.53 22.555 3.53 22.555 1.54 21.16 1.54 21.16 2.43 20.82 2.43  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1
