# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.21 2.27 1.21 2.27 2.16 1.83 2.16  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.015 1.77 1.015 2.39 3.065 2.39 3.065 1.83 4.03 1.83 4.03 3.2 3.69 3.2 3.69 2.09 3.295 2.09 3.295 2.62 0.71 2.62  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.87 1.21 7.21 1.21 7.21 2.16 6.87 2.16  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.72 0.845 11.05 0.845 11.05 4.23 10.72 4.23  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.42 1.595 3.42 1.595 4.59 2.955 4.59 5.225 4.59 5.225 3.42 5.455 3.42 5.455 4.59 7.685 4.59 7.685 3.42 7.915 3.42 7.915 4.59 9.57 4.59 9.57 3.42 9.8 3.42 9.8 4.59 10.37 4.59 11.76 4.59 11.76 5.49 10.37 5.49 2.955 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 9.93 0.45 9.93 1.22 9.7 1.22 9.7 0.45 5.695 0.45 5.695 1.185 5.465 1.185 5.465 0.45 1.595 0.45 1.595 1.185 1.365 1.185 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 2.85 2.955 2.85 2.955 3.19 0.575 3.19 0.575 4.23 0.245 4.23  ;
        POLYGON 3.305 3.42 3.535 3.42 3.535 4 4.26 4 4.26 1.185 3.505 1.185 3.505 0.845 5.235 0.845 5.235 1.415 6.315 1.415 6.315 2.215 6.085 2.215 6.085 1.645 5.005 1.645 5.005 1.075 4.49 1.075 4.49 4.23 3.305 4.23  ;
        POLYGON 4.785 1.875 5.855 1.875 5.855 2.445 6.745 2.445 6.745 2.39 7.605 2.39 7.605 0.845 7.835 0.845 7.835 1.875 9.025 1.875 9.025 2.215 7.835 2.215 7.835 2.62 6.895 2.62 6.895 4.23 6.665 4.23 6.665 2.675 5.625 2.675 5.625 2.215 4.785 2.215  ;
        POLYGON 8.5 2.975 9.255 2.975 9.255 1.79 9.24 1.79 9.24 1.225 8.355 1.225 8.355 0.885 9.47 0.885 9.47 1.705 10.37 1.705 10.37 2.215 10.14 2.215 10.14 1.935 9.485 1.935 9.485 3.205 8.73 3.205 8.73 4.23 8.5 4.23  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_1
