# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__or4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6945 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 1.77 1.015 1.77 1.015 2.555 0.785 2.555 0.785 2.15 0.15 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6945 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.77 2.215 1.77 2.215 2.555 1.83 2.555  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6945 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.95 1.77 3.385 1.77 3.385 2.555 2.95 2.555  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6945 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.07 1.21 4.575 1.21 4.575 2.555 4.345 2.555 4.345 1.59 4.07 1.59  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.285 0.68 6.615 0.68 6.615 4.36 6.285 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 5.265 4.59 5.265 3.79 5.495 3.79 5.495 4.59 5.99 4.59 7.28 4.59 7.28 5.49 5.99 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 5.495 0.45 5.495 0.94 5.265 0.94 5.265 0.45 2.895 0.45 2.895 1.015 2.665 1.015 2.665 0.45 0.475 0.45 0.475 1.015 0.245 1.015 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.29 3.845 4.805 3.845 4.805 0.93 3.84 0.93 3.84 1.475 1.545 1.475 1.545 0.68 1.775 0.68 1.775 1.245 3.61 1.245 3.61 0.7 5.035 0.7 5.035 2.27 5.99 2.27 5.99 2.5 5.035 2.5 5.035 4.075 0.29 4.075  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_1
