* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(((A1 + A2) * (B1 + B2)) * (C1 + C2))
M_i_4_1 net_1 C1 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_5_1 VSS C2 net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_5_0 net_1 C2 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4_0 VSS C1 net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_0 net_1 B1 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_0 net_0 B2 net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_1 net_1 B2 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_1 net_0 B1 net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_10_1 net_4_1 C1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_11_1 VDD C2 net_4_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_11_0 net_4_0 C2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_10_0 ZN C1 net_4_0 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8_0 net_3_1 B1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_0 VDD B2 net_3_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_1 net_3_0 B2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8_1 ZN B1 net_3_0 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_0 net_2_1 A1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_7_0 VDD A2 net_2_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_7_1 net_2_0 A2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_1 ZN A1 net_2_0 VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
