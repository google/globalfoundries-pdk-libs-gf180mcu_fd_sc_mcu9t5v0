# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.16 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.51 2.33 4.55 2.33 4.55 2.71 3.51 2.71  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.15 2.265 14.975 2.265 14.975 2.71 14.15 2.71  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.63 1.77 1.53 1.77 1.53 2.15 0.63 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 18.07 0.845 18.375 0.845 18.375 3.685 18.145 3.685 18.145 1.59 18.07 1.59  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.425 1.495 3.425 1.495 4.59 2.035 4.59 3.005 4.59 3.005 3.905 3.235 3.905 3.235 4.59 7.245 4.59 7.245 3.905 7.475 3.905 7.475 4.59 9.725 4.59 9.725 3.905 9.955 3.905 9.955 4.59 11.535 4.59 13.805 4.59 13.805 3.915 14.035 3.915 14.035 4.59 16.345 4.59 16.345 3.175 16.575 3.175 16.575 4.59 17.07 4.59 17.915 4.59 19.165 4.59 19.165 3.875 19.395 3.875 19.395 4.59 20.16 4.59 20.16 5.49 17.915 5.49 17.07 5.49 11.535 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 20.16 -0.45 20.16 0.45 19.495 0.45 19.495 1.165 19.265 1.165 19.265 0.45 16.535 0.45 16.535 1.42 16.305 1.42 16.305 0.45 7.655 0.45 7.655 1.425 7.425 1.425 7.425 0.45 3.455 0.45 3.455 1.425 3.225 1.425 3.225 0.45 1.595 0.45 1.595 1.08 1.365 1.08 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 2.875 1.805 2.875 1.805 1.54 0.245 1.54 0.245 1.17 0.475 1.17 0.475 1.31 2.035 1.31 2.035 3.105 0.475 3.105 0.475 3.685 0.245 3.685  ;
        POLYGON 3.05 1.87 3.685 1.87 3.685 1.315 4.575 1.315 4.575 1.655 3.915 1.655 3.915 2.1 3.28 2.1 3.28 2.985 4.53 2.985 4.53 3.215 3.05 3.215  ;
        POLYGON 5.265 1.315 5.695 1.315 5.695 1.83 8.19 1.83 8.19 2.06 5.495 2.06 5.495 3.215 5.265 3.215  ;
        POLYGON 6.53 2.47 9.425 2.47 9.425 1.315 9.655 1.315 9.655 2.47 11.095 2.47 11.095 3.215 10.865 3.215 10.865 2.7 8.715 2.7 8.715 3.215 8.485 3.215 8.485 2.7 6.53 2.7  ;
        POLYGON 2.285 1.17 2.715 1.17 2.715 3.445 11.535 3.445 11.535 4.315 11.305 4.315 11.305 3.675 5.99 3.675 5.99 4.26 5.65 4.26 5.65 3.675 2.515 3.675 2.515 3.685 2.285 3.685  ;
        POLYGON 13.085 2.875 13.69 2.875 13.69 1.545 11.845 1.545 11.845 1.205 13.92 1.205 13.92 2.985 15.105 2.985 15.105 2.905 15.335 2.905 15.335 3.245 15.105 3.245 15.105 3.215 13.085 3.215  ;
        POLYGON 10.725 1.315 10.955 1.315 10.955 1.775 12.115 1.775 12.115 3.455 14.225 3.455 14.225 3.475 15.885 3.475 15.885 2.5 17.07 2.5 17.07 2.73 16.115 2.73 16.115 3.705 14.13 3.705 14.13 3.685 11.885 3.685 11.885 2.005 10.725 2.005  ;
        POLYGON 15.685 1.93 17.425 1.93 17.425 1.315 17.655 1.315 17.655 1.975 17.915 1.975 17.915 2.315 17.595 2.315 17.595 3.715 17.365 3.715 17.365 2.27 15.685 2.27  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1
