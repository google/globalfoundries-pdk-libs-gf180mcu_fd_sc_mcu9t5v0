* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__latrsnq_1 D E RN SETN Q VDD VNW VPW VSS
*.PININFO D:I E:I RN:I SETN:I Q:O VDD:P VNW:P VPW:P VSS:G
M_tn3 net8 E VSS VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn9 net2 RN VSS VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn8 net3 D net2 VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn7 net3 E net4 VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn6 net4 net8 net5 VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn5 net6 net1 net5 VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn0 VSS RN net6 VPW nfet_05v0 W=0.700000U L=0.600000U
M_tn11 VSS net4 net0 VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn10 net0 SETN net1 VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn4 net7 net1 VSS VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn1 Q net7 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_tp2 net8 E VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp8 VDD RN net4 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp6 net9 D VDD VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp5 net4 net8 net9 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp4 net10 E net4 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp3 net10 net1 VDD VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp10 VDD net4 net1 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp9 net1 SETN VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp7 net7 net1 VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp0 Q net7 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
