# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.68 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.51 4.455 1.51 4.455 2.025 4.225 2.025 4.225 1.74 2.17 1.74 2.17 2.2 1.83 2.2  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.91 1.915 1.14 1.915 1.14 2.89 3.44 2.89 3.67 2.89 3.67 2.255 5.19 2.255 5.19 1.97 5.53 1.97 5.53 2.485 3.9 2.485 3.9 3.27 3.44 3.27 0.91 3.27  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.09 2.37 9.54 2.37 9.67 2.37 9.67 2.33 10.71 2.33 10.71 2.71 9.54 2.71 8.09 2.71  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.772 ;
    PORT
      LAYER METAL1 ;
        POLYGON 12.845 3.415 13.57 3.415 13.8 3.415 13.8 1.67 12.845 1.67 12.845 0.845 13.29 0.845 13.29 1.44 15.085 1.44 15.085 0.845 15.315 0.845 15.315 3.685 14.985 3.685 14.985 1.67 14.03 1.67 14.03 3.645 13.57 3.645 13.075 3.645 13.075 4.32 12.845 4.32  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.51 2.665 3.51 2.665 4.59 3.44 4.59 6.055 4.59 6.545 4.59 6.545 3.45 6.775 3.45 6.775 4.59 8.815 4.59 8.815 4.35 9.045 4.35 9.045 4.59 12.025 4.59 12.025 4.35 12.255 4.35 12.255 4.59 13.57 4.59 13.865 4.59 13.865 3.875 14.095 3.875 14.095 4.59 15.68 4.59 15.68 5.49 13.57 5.49 6.055 5.49 3.44 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 15.68 -0.45 15.68 0.45 14.195 0.45 14.195 1.165 13.965 1.165 13.965 0.45 8.815 0.45 8.815 1.185 8.585 1.185 8.585 0.45 6.055 0.45 6.055 1.185 5.825 1.185 5.825 0.45 2.715 0.45 2.715 1.185 2.485 1.185 2.485 0.45 0.475 0.45 0.475 1.185 0.245 1.185 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 1.455 1.365 1.455 1.365 0.845 1.6 0.845 1.6 2.43 3.1 2.43 3.1 1.97 3.44 1.97 3.44 2.66 1.37 2.66 1.37 1.685 0.575 1.685 0.575 3.85 0.345 3.85  ;
        POLYGON 3.785 3.51 4.015 3.51 4.015 4.13 5.825 4.13 5.825 3.175 6.055 3.175 6.055 4.36 3.785 4.36  ;
        POLYGON 6.49 0.9 7.795 0.9 7.795 1.91 9.54 1.91 9.54 2.14 7.795 2.14 7.795 3.235 7.565 3.235 7.565 1.13 6.49 1.13  ;
        POLYGON 4.805 2.715 7.005 2.715 7.005 1.645 4.685 1.645 4.685 1.13 3.73 1.13 3.73 0.9 4.915 0.9 4.915 1.415 7.235 1.415 7.235 3.465 10.94 3.465 10.94 2.18 11.73 2.18 11.73 2.41 11.17 2.41 11.17 3.695 7.005 3.695 7.005 2.945 5.035 2.945 5.035 3.9 4.805 3.9  ;
        POLYGON 9.885 0.68 12.355 0.68 12.355 1.49 12.125 1.49 12.125 0.91 10.115 0.91 10.115 1.655 9.885 1.655  ;
        POLYGON 9.93 3.925 11.265 3.925 11.265 3.905 11.71 3.905 11.71 2.64 11.96 2.64 11.96 1.95 11.005 1.95 11.005 1.14 11.235 1.14 11.235 1.72 12.185 1.72 12.185 1.9 13.57 1.9 13.57 2.13 12.19 2.13 12.19 2.87 11.94 2.87 11.94 4.135 11.36 4.135 11.36 4.155 9.93 4.155  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_2
