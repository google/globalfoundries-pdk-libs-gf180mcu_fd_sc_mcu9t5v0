* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__dffsnq_1 D SETN CLK Q VDD VNW VPW VSS
*.PININFO D:I SETN:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G
M_tn3 ncki CLK VSS VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn0 cki ncki VSS VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn10 net13 D VSS VPW nfet_05v0 W=0.590000U L=0.600000U
M_tn6 net13 ncki net3 VPW nfet_05v0 W=0.590000U L=0.600000U
M_tn4 net3 cki net14 VPW nfet_05v0 W=0.590000U L=0.600000U
M_tn5 VSS net4 net14 VPW nfet_05v0 W=0.590000U L=0.600000U
M_tn2 net0 net3 VSS VPW nfet_05v0 W=0.590000U L=0.600000U
M_tn1 net4 SETN net0 VPW nfet_05v0 W=0.590000U L=0.600000U
M_tn13 net5 cki net4 VPW nfet_05v0 W=0.590000U L=0.600000U
M_tn12 net7 ncki net5 VPW nfet_05v0 W=0.590000U L=0.600000U
M_tn14 net1 SETN net7 VPW nfet_05v0 W=0.590000U L=0.600000U
M_tn15 VSS net6 net1 VPW nfet_05v0 W=0.590000U L=0.600000U
M_tn18 net6 net5 VSS VPW nfet_05v0 W=0.750000U L=0.600000U
M_tn16 VSS net6 Q VPW nfet_05v0 W=1.320000U L=0.600000U
M_tp4 ncki CLK VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp0 cki ncki VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp8 VDD D net13 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp9 net3 cki net13 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp6 net10 ncki net3 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net10 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp3 net4 net3 VDD VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp2 VDD SETN net4 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp18 net5 ncki net4 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp17 net7 cki net5 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp12 net7 SETN VDD VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp13 VDD net6 net7 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp16 net6 net5 VDD VNW pfet_05v0 W=1.100000U L=0.500000U
M_tp14 VDD net6 Q VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
