* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__dlya_2 I Z VDD VNW VPW VSS
*.PININFO I:I Z:O VDD:P VNW:P VPW:P VSS:G
*.EQN Z=I
M_i_2_0 Z_neg I VSS VPW nfet_05v0 W=0.360000U L=0.600000U
M_i_2 VSS Z_neg net_2 VPW nfet_05v0 W=0.360000U L=0.600000U
M_i_3_6 net_3 net_2 VSS VPW nfet_05v0 W=0.360000U L=0.600000U
M_i_2_0_18 Z net_3 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_0_18_1 Z net_3 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_0 Z_neg I VDD VNW pfet_05v0 W=0.360000U L=0.500000U
M_i_1 VDD Z_neg net_2 VNW pfet_05v0 W=0.360000U L=0.500000U
M_i_0_29 net_3 net_2 VDD VNW pfet_05v0 W=0.360000U L=0.500000U
M_i_3_0_0 Z net_3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_3_0_0_14 Z net_3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
