# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 24.64 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.055 2.33 3.89 2.33 3.89 2.71 3.055 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.95 2.48 17.515 2.48 17.515 2.71 17.21 2.71 17.21 3.27 16.95 3.27  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.27 1.77 15.53 1.77 15.53 2.765 15.27 2.765  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.295 1.57 2.295 1.57 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.59 2.875 22.435 2.875 22.665 2.875 22.665 1.655 20.59 1.655 20.59 0.845 20.82 0.845 20.82 1.395 22.55 1.395 22.55 0.815 23.06 0.815 23.06 3.685 22.63 3.685 22.63 3.105 22.435 3.105 20.82 3.105 20.82 3.685 20.59 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.205 4.59 3.205 3.515 3.435 3.515 3.435 4.59 7.465 4.59 7.465 4.49 7.695 4.49 7.695 4.59 10.665 4.59 10.665 4.49 10.895 4.49 10.895 4.59 12.63 4.59 14.695 4.59 14.695 3.96 15.035 3.96 15.035 4.59 16.735 4.59 16.735 3.96 17.075 3.96 17.075 4.59 18.5 4.59 18.83 4.59 18.83 3.435 19.06 3.435 19.06 4.59 19.57 4.59 19.57 3.875 19.8 3.875 19.8 4.59 21.61 4.59 21.61 3.875 21.84 3.875 21.84 4.59 22.435 4.59 23.65 4.59 23.65 3.875 23.88 3.875 23.88 4.59 24.64 4.59 24.64 5.49 22.435 5.49 18.5 5.49 12.63 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 24.64 -0.45 24.64 0.45 24.18 0.45 24.18 1.165 23.95 1.165 23.95 0.45 21.94 0.45 21.94 1.165 21.71 1.165 21.71 0.45 19.7 0.45 19.7 1.165 19.47 1.165 19.47 0.45 17.02 0.45 17.02 1.225 16.79 1.225 16.79 0.45 8.635 0.45 8.635 1.425 8.405 1.425 8.405 0.45 3.435 0.45 3.435 1.425 3.205 1.425 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.225 1.315 4.555 1.315 4.555 3.685 4.225 3.685  ;
        POLYGON 6.285 3.35 8.935 3.35 8.935 3.8 6.285 3.8  ;
        POLYGON 5.245 1.315 5.675 1.315 5.675 2.685 9.865 2.685 9.865 2.575 10.095 2.575 10.095 2.915 5.475 2.915 5.475 3.685 5.245 3.685  ;
        POLYGON 9.425 3.46 11.285 3.46 11.285 2.345 7.095 2.345 7.095 2.455 6.865 2.455 6.865 2.115 11.285 2.115 11.285 1.315 11.515 1.315 11.515 3.57 11.905 3.57 11.905 2.875 12.135 2.875 12.135 3.8 9.425 3.8  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 3.055 3.895 3.055 3.895 4.03 12.63 4.03 12.63 4.26 3.665 4.26 3.665 3.285 2.615 3.285 2.615 3.685 2.385 3.685  ;
        POLYGON 6.125 1.655 10.825 1.655 10.825 0.68 14.455 0.68 14.455 0.91 11.055 0.91 11.055 1.885 6.355 1.885 6.355 2.115 6.125 2.115  ;
        POLYGON 13.525 1.31 16 1.31 16 3.225 15.77 3.225 15.77 1.54 14.175 1.54 14.175 3.215 13.945 3.215 13.945 1.655 13.525 1.655  ;
        POLYGON 12.405 1.315 13.155 1.315 13.155 3.5 18.27 3.5 18.27 2.425 18.5 2.425 18.5 3.73 12.925 3.73 12.925 1.655 12.405 1.655  ;
        POLYGON 16.295 1.83 18.75 1.83 18.75 1.315 18.98 1.315 18.98 1.775 20.24 1.775 20.24 2.005 22.435 2.005 22.435 2.29 20.01 2.29 20.01 2.115 18.04 2.115 18.04 3.225 17.81 3.225 17.81 2.06 16.295 2.06  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4
