# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai33_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai33_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.59 2.28 9.93 2.28 9.93 2.71 9.59 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.55 1.77 8.81 1.77 8.81 1.82 10.39 1.82 10.39 2.27 12.22 2.27 12.22 2.5 10.16 2.5 10.16 2.05 8.89 2.05 8.89 2.5 8.55 2.5  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 2.215 7.735 2.215 7.735 2.94 13.005 2.94 13.005 2.215 13.235 2.215 13.235 3.17 7.43 3.17  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 2.27 3.26 2.27 3.26 2.71 2.92 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.99 2.27 2.39 2.27 2.39 1.77 3.72 1.77 3.72 2.27 5.5 2.27 5.5 2.5 3.49 2.5 3.49 2 2.65 2 2.65 2.5 1.99 2.5  ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.94 5.73 2.94 5.73 2.27 6.62 2.27 6.62 2.5 5.96 2.5 5.96 3.17 0.71 3.17  ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.3284 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.655 3.4 13.465 3.4 13.465 1.59 10.23 1.59 10.23 1.48 8.03 1.48 8.03 1.25 10.23 1.25 10.23 1.14 10.555 1.14 10.555 1.25 13.695 1.25 13.695 3.63 10.505 3.63 10.505 4.36 10.275 4.36 10.275 3.63 3.885 3.63 3.885 4.36 3.655 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.86 0.575 3.86 0.575 4.59 6.915 4.59 6.915 3.86 7.145 3.86 7.145 4.59 13.585 4.59 13.585 3.86 13.815 3.86 13.815 4.59 13.915 4.59 14.56 4.59 14.56 5.49 13.915 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 6.075 0.45 6.075 1.565 5.845 1.565 5.845 0.45 3.835 0.45 3.835 1 3.605 1 3.605 0.45 1.595 0.45 1.595 1.455 1.365 1.455 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 1.685 1.93 1.685 1.93 0.73 2.715 0.73 2.715 1.31 4.725 1.31 4.725 0.73 4.955 0.73 4.955 1.795 6.965 1.795 6.965 0.68 13.915 0.68 13.915 1.02 11.445 1.02 11.445 0.91 9.435 0.91 9.435 1.02 7.195 1.02 7.195 2.025 4.725 2.025 4.725 1.54 2.16 1.54 2.16 1.915 0.245 1.915  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai33_2
