# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.36 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.67 1.755 12.595 1.755 12.595 2.27 14.23 2.27 14.23 2.5 12.365 2.5 12.365 1.985 10.15 1.985 10.15 2.5 9.67 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.93 2.27 9.27 2.27 9.27 2.73 11.35 2.73 11.35 2.215 12.135 2.215 12.135 2.73 15.705 2.73 15.705 2.215 15.935 2.215 15.935 2.96 8.93 2.96  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.27 1.05 2.27 1.05 2.73 3.745 2.73 3.745 2.215 3.975 2.215 3.975 2.73 6.3 2.73 6.3 2.27 8.11 2.27 8.11 2.5 6.53 2.5 6.53 2.96 0.71 2.96  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.728 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.755 4.435 1.755 4.435 2.27 6.07 2.27 6.07 2.5 4.205 2.5 4.205 1.985 2.17 1.985 2.17 2.5 1.83 2.5  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.6976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 3.19 16.165 3.19 16.165 1.425 10.39 1.425 10.39 1.195 16.395 1.195 16.395 3.42 15.775 3.42 15.775 4.36 15.545 4.36 15.545 3.42 13.735 3.42 13.735 4.36 13.505 4.36 13.505 3.42 11.695 3.42 11.695 4.36 11.465 4.36 11.465 3.42 9.655 3.42 9.655 4.36 9.425 4.36 9.425 3.42 7.615 3.42 7.615 4.36 7.385 4.36 7.385 3.42 5.575 3.42 5.575 4.36 5.345 4.36 5.345 3.42 3.535 3.42 3.535 4.36 2.89 4.36 2.89 3.42 1.495 3.42 1.495 4.36 1.265 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.65 0.475 3.65 0.475 4.59 2.285 4.59 2.285 3.65 2.515 3.65 2.515 4.59 4.325 4.59 4.325 3.65 4.555 3.65 4.555 4.59 6.365 4.59 6.365 3.65 6.595 3.65 6.595 4.59 8.405 4.59 8.405 3.65 8.635 3.65 8.635 4.59 10.445 4.59 10.445 3.65 10.675 3.65 10.675 4.59 12.485 4.59 12.485 3.65 12.715 3.65 12.715 4.59 14.525 4.59 14.525 3.65 14.755 3.65 14.755 4.59 16.565 4.59 16.565 3.65 16.795 3.65 16.795 4.59 16.85 4.59 17.36 4.59 17.36 5.49 16.85 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.36 -0.45 17.36 0.45 6.595 0.45 6.595 1.02 6.365 1.02 6.365 0.45 2.515 0.45 2.515 1.02 2.285 1.02 2.285 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 1.26 4.325 1.26 4.325 0.68 4.555 0.68 4.555 1.26 9.93 1.26 9.93 0.735 16.85 0.735 16.85 0.965 10.16 0.965 10.16 1.49 0.245 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nand4_4
