# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.4 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.87 2.27 7.29 2.27 7.29 2.71 6.87 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.75 2.27 6.18 2.27 6.18 2.71 5.75 2.71  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.51 1.77 3.98 1.77 3.98 2.5 3.51 2.5  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.63 2.27 5.05 2.27 5.05 2.71 4.63 2.71  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 2.15 2.09 2.15 2.09 2.71 1.83 2.71  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.71 0.71 2.71  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.9438 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.64 3.55 7.815 3.55 7.815 4.36 7.585 4.36 7.585 3.83 4.555 3.83 3.485 3.83 3.485 4.36 3.255 4.36 3.255 3.45 4.555 3.45 6.41 3.45 6.41 1.14 6.795 1.14 6.795 1.48 6.64 1.48  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 4.555 4.59 5.345 4.59 5.345 4.06 5.575 4.06 5.575 4.59 7.915 4.59 8.4 4.59 8.4 5.49 7.915 5.49 4.555 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 8.4 -0.45 8.4 0.45 2.715 0.45 2.715 1.205 2.485 1.205 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.365 0.68 1.595 0.68 1.595 1.435 3.1 1.435 3.1 1.31 4.325 1.31 4.325 1.14 4.555 1.14 4.555 1.54 3.305 1.54 3.305 1.665 1.365 1.665  ;
        POLYGON 3.15 0.68 7.915 0.68 7.915 1.49 7.685 1.49 7.685 0.91 5.675 0.91 5.675 1.49 5.445 1.49 5.445 0.91 3.49 0.91 3.49 0.965 3.15 0.965  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_1
