# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.68 BY 5.04 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.625 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.23 1.21 10.425 1.21 10.49 1.21 10.49 2.405 10.425 2.405 10.23 2.405  ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.21 1.77 2.09 1.77 2.09 2.35 1.21 2.35  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.4716 ;
    PORT
      LAYER METAL1 ;
        POLYGON 13.59 2.89 13.94 2.89 13.94 1.59 13.59 1.59 13.59 1.21 13.94 1.21 13.94 0.79 14.2 0.79 14.2 3.685 13.59 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.95 4.59 13.49 4.59 15.68 4.59 15.68 5.49 13.49 5.49 2.715 5.49 0 5.49 0 4.59 0.695 4.59 0.695 3.44 0.925 3.44 0.925 4.59 2.715 4.59 5.805 4.59 5.805 3.85 6.035 3.85 6.035 4.59 8.72 4.59 8.72 3.85 11.14 3.85 11.14 4.02 12.95 4.02 12.95 3.44 13.18 3.44 13.18 4.02 13.49 4.02 14.99 4.02 14.99 3.44 15.22 3.44 15.22 4.25 13.49 4.25 8.95 4.25  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 15.68 -0.45 15.68 0.45 15.29 0.45 15.29 1.43 15.06 1.43 15.06 0.45 13.05 0.45 13.05 1.43 12.82 1.43 12.82 0.45 9.25 0.45 9.25 1.13 9.02 1.13 9.02 0.45 5.85 0.45 5.85 1.13 5.62 1.13 5.62 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.79 0.475 0.79 0.475 1.305 2.485 1.305 2.485 0.79 2.715 0.79 2.715 1.535 0.245 1.535  ;
        POLYGON 3.445 1.79 3.675 1.79 3.675 2.485 4.77 2.485 4.77 2.715 3.445 2.715  ;
        POLYGON 3.215 2.945 5 2.945 5 1.605 6.345 1.605 6.345 2.35 6.005 2.35 6.005 1.835 5.23 1.835 5.23 3.175 3.785 3.175 3.785 4.25 3.555 4.25 3.555 3.175 2.985 3.175 2.985 0.845 3.89 0.845 3.89 1.075 3.215 1.075  ;
        POLYGON 7.4 0.845 8.185 0.845 8.185 1.075 7.63 1.075 7.63 2.93 7.985 2.93 7.985 3.16 7.4 3.16  ;
        POLYGON 8.225 2.12 9.685 2.12 9.685 0.75 10.425 0.75 10.425 0.98 9.915 0.98 9.915 2.93 10.025 2.93 10.025 3.16 9.685 3.16 9.685 2.35 8.225 2.35  ;
        POLYGON 5.46 2.065 5.69 2.065 5.69 3.39 6.74 3.39 6.74 0.79 6.97 0.79 6.97 3.39 11.47 3.39 11.47 2.12 12.425 2.12 12.425 2.35 11.7 2.35 11.7 3.62 7.055 3.62 7.055 4.25 6.825 4.25 6.825 3.62 5.46 3.62  ;
        POLYGON 11.93 2.875 12.655 2.875 12.655 1.89 10.86 1.89 10.86 0.79 11.09 0.79 11.09 1.66 12.885 1.66 12.885 2.065 13.49 2.065 13.49 2.405 12.885 2.405 12.885 3.105 12.16 3.105 12.16 3.685 11.93 3.685  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_2
