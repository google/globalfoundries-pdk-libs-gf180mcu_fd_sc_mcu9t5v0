* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1 D RN SETN CLKN Q VDD VNW VPW VSS
*.PININFO D:I RN:I SETN:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G
M_tn2 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn1 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn0 net14 D VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net14 cki net3 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net3 ncki net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net15 net4 net16 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS RN net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 net0 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net4 SETN net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net5 ncki net4 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn13 net7 cki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net1 SETN net7 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 VSS net6 net1 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn18 net2 RN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn17 net6 net5 net2 VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn19 Q net6 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp2 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp1 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp0 VDD D net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net3 ncki net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net13 cki net3 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 VDD net4 net13 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net13 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp4 VDD net3 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 VDD SETN net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp20 net4 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp19 net5 ncki net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net7 SETN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp14 net7 net6 VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp16 net6 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 VDD net5 net6 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp17 Q net6 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
