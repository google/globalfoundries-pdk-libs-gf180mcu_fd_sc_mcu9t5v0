# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__hold
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__hold 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.04 BY 5.04 ;
  PIN Z
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.4896 ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 1.415 3.95 1.415 3.95 2.575 3.51 2.575 3.51 1.645 0.575 1.645 0.575 3.605 0.245 3.605  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 3.225 4.59 3.225 3.265 3.455 3.265 3.455 4.59 4.575 4.59 5.04 4.59 5.04 5.49 4.575 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.04 -0.45 5.04 0.45 3.455 0.45 3.455 1.185 3.225 1.185 3.225 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.51 1.875 2.85 1.875 2.85 2.805 4.345 2.805 4.345 0.845 4.575 0.845 4.575 4.075 4.245 4.075 4.245 3.035 2.51 3.035  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__hold
