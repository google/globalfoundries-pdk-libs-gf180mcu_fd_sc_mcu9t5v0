# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtp_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtp_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.625 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.23 1.77 10.315 1.77 10.49 1.77 10.49 2.71 10.315 2.71 10.23 2.71  ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.175 2.09 2.175 2.09 2.405 0.97 2.405 0.97 2.71 0.71 2.71  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.415 1.77 0.415 2.71 0.15 2.71  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.9432 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.885 2.875 15.37 2.875 15.955 2.875 15.955 1.745 13.885 1.745 13.885 0.795 14.115 0.795 14.115 1.515 15.77 1.515 15.77 0.71 16.355 0.71 16.355 3.685 15.955 3.685 15.955 3.105 15.37 3.105 14.145 3.105 14.145 3.685 13.885 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.125 4.59 15.37 4.59 17.92 4.59 17.92 5.49 15.37 5.49 2.715 5.49 0 5.49 0 4.59 0.625 4.59 0.625 3.44 0.855 3.44 0.855 4.59 2.715 4.59 5.805 4.59 5.805 3.855 6.035 3.855 6.035 4.59 8.865 4.59 8.865 3.855 9.095 3.855 9.095 4.59 10.855 4.59 10.855 3.855 11.085 3.855 11.085 4.59 12.895 4.59 12.895 3.44 13.125 3.44 13.125 4.02 14.935 4.02 14.935 3.44 15.165 3.44 15.165 4.02 15.37 4.02 16.975 4.02 16.975 3.44 17.205 3.44 17.205 4.25 15.37 4.25 13.125 4.25  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 17.475 0.45 17.475 1.485 17.245 1.485 17.245 0.45 15.235 0.45 15.235 1.035 15.005 1.035 15.005 0.45 12.995 0.45 12.995 1.485 12.765 1.485 12.765 0.45 9.195 0.45 9.195 1.135 8.965 1.135 8.965 0.45 5.795 0.45 5.795 1.135 5.565 1.135 5.565 0.45 1.65 0.45 1.65 1.08 1.31 1.08 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.795 0.475 0.795 0.475 1.31 2.485 1.31 2.485 0.795 2.715 0.795 2.715 1.54 0.245 1.54  ;
        POLYGON 3.445 1.79 4.715 1.79 4.715 2.77 4.485 2.77 4.485 2.13 3.445 2.13  ;
        POLYGON 3.215 2.82 4.26 2.82 4.26 3 4.945 3 4.945 1.66 6.095 1.66 6.095 2.175 6.53 2.175 6.53 2.405 5.865 2.405 5.865 1.89 5.175 1.89 5.175 3.23 4.265 3.23 4.265 4.25 4.035 4.25 4.035 3.05 2.985 3.05 2.985 0.85 3.89 0.85 3.89 1.08 3.215 1.08  ;
        POLYGON 7.345 2.12 7.845 2.12 7.845 0.795 8.13 0.795 8.13 3.16 7.79 3.16 7.79 2.46 7.345 2.46  ;
        POLYGON 8.37 2.175 9.77 2.175 9.77 1.31 10.085 1.31 10.085 0.795 10.315 0.795 10.315 1.54 10 1.54 10 2.935 10.17 2.935 10.17 3.165 9.77 3.165 9.77 2.405 8.37 2.405  ;
        POLYGON 5.405 2.12 5.635 2.12 5.635 3.395 6.76 3.395 6.76 1.135 6.685 1.135 6.685 0.795 6.99 0.795 6.99 3.395 11.415 3.395 11.415 2.175 12.6 2.175 12.6 2.405 11.645 2.405 11.645 3.625 7.055 3.625 7.055 4.25 6.825 4.25 6.825 3.625 5.405 3.625  ;
        POLYGON 11.875 2.875 12.83 2.875 12.83 1.945 10.805 1.945 10.805 0.795 11.035 0.795 11.035 1.715 13.06 1.715 13.06 1.975 15.37 1.975 15.37 2.315 13.06 2.315 13.06 3.105 12.105 3.105 12.105 3.685 11.875 3.685  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtp_4
