# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 34.72 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.53 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.685 2.215 9.845 2.215 9.845 2.65 0.685 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 15.506 ;
    PORT
      LAYER METAL1 ;
        POLYGON 12.745 3.09 21.225 3.09 22.465 3.09 22.465 1.745 12.745 1.745 12.745 0.945 13.005 0.945 13.005 1.515 14.985 1.515 14.985 0.945 15.215 0.945 15.215 1.515 17.225 1.515 17.225 0.945 17.455 0.945 17.455 1.515 19.465 1.515 19.465 0.945 19.695 0.945 19.695 1.515 21.705 1.515 21.705 0.945 21.935 0.945 21.935 1.445 23.945 1.445 23.945 0.945 24.175 0.945 24.175 1.445 26.185 1.445 26.185 0.945 26.415 0.945 26.415 1.445 28.425 1.445 28.425 0.945 28.655 0.945 28.655 1.445 30.665 1.445 30.665 0.945 30.895 0.945 30.895 1.445 32.905 1.445 32.905 0.945 33.135 0.945 33.135 1.675 23.215 1.675 23.215 3.09 32.605 3.09 33.035 3.09 33.035 4.36 32.805 4.36 32.805 3.32 32.605 3.32 30.795 3.32 30.795 4.36 30.565 4.36 30.565 3.32 28.555 3.32 28.555 4.36 28.325 4.36 28.325 3.32 26.315 3.32 26.315 4.36 26.085 4.36 26.085 3.32 24.075 3.32 24.075 4.36 23.845 4.36 23.845 3.32 21.835 3.32 21.835 4.36 21.605 4.36 21.605 3.32 21.225 3.32 19.595 3.32 19.595 4.36 19.365 4.36 19.365 3.32 17.355 3.32 17.355 4.36 17.125 4.36 17.125 3.32 15.115 3.32 15.115 4.36 14.885 4.36 14.885 3.32 12.975 3.32 12.975 4.36 12.745 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.875 11.575 3.875 11.575 4.59 13.765 4.59 13.765 3.55 13.995 3.55 13.995 4.59 16.005 4.59 16.005 3.55 16.235 3.55 16.235 4.59 18.245 4.59 18.245 3.55 18.475 3.55 18.475 4.59 20.485 4.59 20.485 3.55 20.715 3.55 20.715 4.59 21.225 4.59 22.725 4.59 22.725 3.55 22.955 3.55 22.955 4.59 24.965 4.59 24.965 3.55 25.195 3.55 25.195 4.59 27.205 4.59 27.205 3.55 27.435 3.55 27.435 4.59 29.445 4.59 29.445 3.55 29.675 3.55 29.675 4.59 31.685 4.59 31.685 3.55 31.915 3.55 31.915 4.59 32.605 4.59 33.925 4.59 33.925 3.55 34.155 3.55 34.155 4.59 34.72 4.59 34.72 5.49 32.605 5.49 21.225 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 34.72 -0.45 34.72 0.45 34.255 0.45 34.255 1.285 34.025 1.285 34.025 0.45 32.015 0.45 32.015 1.215 31.785 1.215 31.785 0.45 29.775 0.45 29.775 1.215 29.545 1.215 29.545 0.45 27.535 0.45 27.535 1.215 27.305 1.215 27.305 0.45 25.295 0.45 25.295 1.215 25.065 1.215 25.065 0.45 23.055 0.45 23.055 1.215 22.825 1.215 22.825 0.45 20.815 0.45 20.815 1.215 20.585 1.215 20.585 0.45 18.575 0.45 18.575 1.285 18.345 1.285 18.345 0.45 16.335 0.45 16.335 1.285 16.105 1.285 16.105 0.45 14.095 0.45 14.095 1.285 13.865 1.285 13.865 0.45 11.675 0.45 11.675 1.285 11.445 1.285 11.445 0.45 9.435 0.45 9.435 1.285 9.205 1.285 9.205 0.45 7.195 0.45 7.195 1.285 6.965 1.285 6.965 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.365 3.09 10.225 3.09 10.225 1.745 1.365 1.745 1.365 0.945 1.595 0.945 1.595 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 5.845 1.515 5.845 0.945 6.075 0.945 6.075 1.515 8.085 1.515 8.085 0.945 8.315 0.945 8.315 1.515 10.325 1.515 10.325 0.945 10.555 0.945 10.555 2.215 21.225 2.215 21.225 2.65 10.455 2.65 10.455 4.36 10.225 4.36 10.225 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
        POLYGON 23.445 2.215 32.605 2.215 32.605 2.65 23.445 2.65  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_20
