# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__fill_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fill_32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 17.92 4.59 17.92 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__fill_32
