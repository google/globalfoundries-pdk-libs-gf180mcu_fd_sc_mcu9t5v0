# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.26 1.77 3.26 2.71 2.95 2.71  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.895 1.835 1.37 1.835 1.37 1.31 4.07 1.31 4.07 1.21 4.33 1.21 4.33 1.78 5 1.78 5 2.765 5.38 2.765 5.38 2.995 4.77 2.995 4.77 2.15 4.07 2.15 4.07 1.54 1.6 1.54 1.6 2.065 0.895 2.065  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.34 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.475 1.77 2.475 2.065 2.09 2.065 2.09 2.71 1.83 2.71  ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.355 0.845 12.73 0.845 12.73 4.36 12.355 4.36  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.39 4.59 1.39 3.55 1.62 3.55 1.62 4.59 3.13 4.59 3.13 3.86 3.36 3.86 3.36 4.59 6.65 4.59 6.65 3.69 6.88 3.69 6.88 4.59 9.42 4.59 9.42 3.55 9.65 3.55 9.65 4.59 10.04 4.59 11.335 4.59 11.335 3.88 11.565 3.88 11.565 4.59 12.01 4.59 13.375 4.59 13.375 3.88 13.605 3.88 13.605 4.59 14 4.59 14 5.49 12.01 5.49 10.04 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14 -0.45 14 0.45 13.755 0.45 13.755 1.605 13.525 1.605 13.525 0.45 11.515 0.45 11.515 1.605 11.285 1.605 11.285 0.45 9.6 0.45 9.6 1.135 9.37 1.135 9.37 0.45 7.58 0.45 7.58 1.135 7.35 1.135 7.35 0.45 1.775 0.45 1.775 1.08 1.435 1.08 1.435 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.37 0.795 0.6 0.795 0.6 2.94 4.31 2.94 4.31 2.38 4.54 2.38 4.54 3.17 0.6 3.17 0.6 4.36 0.37 4.36  ;
        POLYGON 2.11 3.4 5.12 3.4 5.12 3.8 5.61 3.8 5.61 1.135 4.55 1.135 4.55 0.795 6.67 0.795 6.67 1.365 7.98 1.365 7.98 2.12 7.75 2.12 7.75 1.595 6.44 1.595 6.44 1.025 5.84 1.025 5.84 4.03 4.89 4.03 4.89 3.63 2.34 3.63 2.34 4.03 2.11 4.03  ;
        POLYGON 6.07 1.78 6.3 1.78 6.3 1.89 7.52 1.89 7.52 2.35 8.21 2.35 8.21 0.795 8.88 0.795 8.88 1.78 10.04 1.78 10.04 2.12 8.44 2.12 8.44 4.36 7.895 4.36 7.895 2.58 7.29 2.58 7.29 2.12 6.07 2.12  ;
        POLYGON 10.44 1.225 10.72 1.225 10.72 1.835 12.01 1.835 12.01 2.065 10.67 2.065 10.67 4.36 10.44 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_2
