# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 27.44 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.77 4.33 1.77 4.33 2.215 3.51 2.215  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.97 1.77 0.97 2.215 0.15 2.215  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.07 1.77 18.89 1.77 18.89 2.215 18.07 2.215  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 1.77 2.09 1.77 2.09 2.215 1.27 2.215  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 2.33 6.91 2.33 6.91 2.71 5.75 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.55965 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.59 0.845 23.82 0.845 23.82 1.21 25.83 1.21 25.83 0.845 26.06 0.845 26.06 1.655 23.93 1.655 23.93 2.88 25.92 2.88 25.92 3.69 25.69 3.69 25.69 3.11 23.87 3.11 23.87 3.69 23.59 3.69  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 3.23 1.545 3.23 1.545 4.59 5.085 4.59 5.085 3.4 5.315 3.4 5.315 4.59 7.2 4.59 7.2 4.125 7.54 4.125 7.54 4.59 9.275 4.59 9.72 4.59 12.045 4.59 12.045 4.51 12.275 4.51 12.275 4.59 14.305 4.59 14.305 4.07 14.535 4.07 14.535 4.59 16.235 4.59 18.305 4.59 18.305 3.075 18.535 3.075 18.535 4.59 19.555 4.59 20.565 4.59 20.565 3.88 20.795 3.88 20.795 4.59 22.605 4.59 22.605 3.88 22.835 3.88 22.835 4.59 23.275 4.59 24.66 4.59 24.66 3.88 24.89 3.88 24.89 4.59 26.85 4.59 26.85 3.88 27.08 3.88 27.08 4.59 27.44 4.59 27.44 5.49 23.275 5.49 19.555 5.49 16.235 5.49 9.72 5.49 9.275 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 27.44 -0.45 27.44 0.45 27.18 0.45 27.18 1.655 26.95 1.655 26.95 0.45 24.94 0.45 24.94 0.98 24.71 0.98 24.71 0.45 22.7 0.45 22.7 1.655 22.47 1.655 22.47 0.45 20.46 0.45 20.46 1.265 20.23 1.265 20.23 0.45 12.455 0.45 12.455 1.12 12.225 1.12 12.225 0.45 7.535 0.45 7.535 1.18 7.305 1.18 7.305 0.45 5.735 0.45 5.735 0.53 5.505 0.53 5.505 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.295 2.455 2.545 2.455 2.545 1.54 0.245 1.54 0.245 0.925 0.475 0.925 0.475 1.31 2.775 1.31 2.775 2.455 4.605 2.455 4.605 1.93 4.835 1.93 4.835 2.685 0.525 2.685 0.525 4.04 0.295 4.04  ;
        POLYGON 6.235 3.095 7.14 3.095 7.14 2.1 6.185 2.1 6.185 1.27 6.415 1.27 6.415 1.87 7.98 1.87 7.98 2.215 7.37 2.215 7.37 3.435 6.235 3.435  ;
        POLYGON 3.325 2.94 5.775 2.94 5.775 3.665 9.045 3.665 9.045 3.065 9.275 3.065 9.275 3.895 5.545 3.895 5.545 3.17 3.555 3.17 3.555 4.04 3.325 4.04  ;
        POLYGON 3.325 0.76 6.875 0.76 6.875 1.41 7.965 1.41 7.965 0.76 9.375 0.76 9.375 1.12 9.145 1.12 9.145 0.99 8.195 0.99 8.195 1.64 6.645 1.64 6.645 0.99 3.555 0.99 3.555 1.13 3.325 1.13  ;
        POLYGON 8.275 3.095 8.425 3.095 8.425 1.22 8.655 1.22 8.655 1.985 9.72 1.985 9.72 2.215 8.655 2.215 8.655 3.435 8.275 3.435  ;
        POLYGON 10.065 0.925 10.495 0.925 10.495 1.985 13.17 1.985 13.17 2.215 10.295 2.215 10.295 3.875 10.065 3.875  ;
        POLYGON 10.79 1.525 12.685 1.525 12.685 0.68 15.13 0.68 15.13 0.91 12.915 0.91 12.915 1.755 10.79 1.755  ;
        POLYGON 11.33 2.445 14.405 2.445 14.405 1.315 14.635 1.315 14.635 2.445 15.775 2.445 15.775 3.38 15.545 3.38 15.545 2.675 13.515 2.675 13.515 3.77 13.285 3.77 13.285 2.675 11.33 2.675  ;
        POLYGON 10.59 4.05 13.745 4.05 13.745 3.095 13.975 3.095 13.975 3.61 16.005 3.61 16.005 3.095 16.235 3.095 16.235 4.36 16.005 4.36 16.005 3.84 13.975 3.84 13.975 4.28 10.59 4.28  ;
        POLYGON 17.815 2.615 19.555 2.615 19.555 3.715 19.325 3.715 19.325 2.845 17.815 2.845 17.815 3.9 17.585 3.9 17.585 1.5 16.645 1.5 16.645 1.16 18.32 1.16 18.32 1.5 17.815 1.5  ;
        POLYGON 15.525 1.085 16.185 1.085 16.185 0.7 19.35 0.7 19.35 1.985 21.055 1.985 21.055 2.215 19.12 2.215 19.12 0.93 16.415 0.93 16.415 1.73 16.795 1.73 16.795 3.9 16.565 3.9 16.565 1.96 16.185 1.96 16.185 1.425 15.525 1.425  ;
        POLYGON 19.905 2.445 21.35 2.445 21.35 0.845 21.58 0.845 21.58 2.42 23.275 2.42 23.275 2.76 21.815 2.76 21.815 3.69 21.585 3.69 21.585 2.785 19.905 2.785  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4
