* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I B1:I B2:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(((A1 + A2) * (B1 + B2)) * C)
M_i_3_3 net_1 B1 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4_3 VSS B2 net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4_2 net_1 B2 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_2 VSS B1 net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_1 net_1 B1 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4_1 VSS B2 net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4_0 net_1 B2 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_0 VSS B1 net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_3 net_1 C net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_2 net_0 C net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_1 net_1 C net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_0 net_0 C net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_3 ZN A1 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_3 net_0 A2 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_2 ZN A2 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_2 net_0 A1 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_1 net_0 A2 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_0 ZN A2 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0 net_0 A1 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_8_3 net_3_0 B1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_3 VDD B2 net_3_0 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_2 net_3_1 B2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8_2 ZN B1 net_3_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8_1 net_3_2 B1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_1 VDD B2 net_3_2 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_0 net_3_3 B2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8_0 ZN B1 net_3_3 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_7_3 VDD C ZN VNW pfet_05v0 W=1.460000U L=0.500000U
M_i_7_2 ZN C VDD VNW pfet_05v0 W=1.460000U L=0.500000U
M_i_7_1 VDD C ZN VNW pfet_05v0 W=1.460000U L=0.500000U
M_i_7_0 ZN C VDD VNW pfet_05v0 W=1.460000U L=0.500000U
M_i_5_3 net_2_0 A1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_3 VDD A2 net_2_0 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_2 net_2_1 A2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_5_2 ZN A1 net_2_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_5_1 net_2_2 A1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_1 VDD A2 net_2_2 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_0 net_2_3 A2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_5_0 ZN A1 net_2_3 VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
