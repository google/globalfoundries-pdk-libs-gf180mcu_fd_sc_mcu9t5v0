# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__or4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.035 2.215 4.33 2.215 4.33 2.71 4.035 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.06 2.27 3.67 2.27 3.67 2.94 4.63 2.94 4.63 2.215 6.565 2.215 6.565 2.71 4.86 2.71 4.86 3.17 3.44 3.17 3.44 2.5 3.06 2.5  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 1.755 7.13 1.755 7.13 2.27 7.74 2.27 7.74 2.5 6.87 2.5 6.87 1.985 2.28 1.985 2.28 2.5 1.94 2.5  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.27 1.21 2.27 1.21 2.89 3.21 2.89 3.21 3.4 7.97 3.4 7.97 2.27 8.86 2.27 8.86 2.5 8.2 2.5 8.2 3.63 0.87 3.63  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.5505 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.17 3.295 11.05 3.295 11.28 3.295 11.28 1.95 10.505 1.95 10.505 0.68 10.735 0.68 10.735 1.72 12.745 1.72 12.745 0.68 12.975 0.68 12.975 1.95 11.835 1.95 11.835 3.295 12.875 3.295 12.875 4.36 12.645 4.36 12.645 3.525 11.05 3.525 10.735 3.525 10.735 4.36 10.17 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.755 0.575 3.755 0.575 4.59 9.46 4.59 9.46 4.275 9.69 4.275 9.69 4.59 11.05 4.59 11.575 4.59 11.575 3.755 11.805 3.755 11.805 4.59 13.765 4.59 13.765 3.755 13.995 3.755 13.995 4.59 14.56 4.59 14.56 5.49 11.05 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 14.095 0.45 14.095 1.49 13.865 1.49 13.865 0.45 11.855 0.45 11.855 1.49 11.625 1.49 11.625 0.45 9.435 0.45 9.435 1.02 9.205 1.02 9.205 0.45 7.195 0.45 7.195 1.02 6.965 1.02 6.965 0.45 4.955 0.45 4.955 1.02 4.725 1.02 4.725 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.02 0.245 1.02 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 4.72 3.86 9.09 3.86 9.09 1.48 1.365 1.48 1.365 0.68 1.595 0.68 1.595 1.25 3.605 1.25 3.605 0.68 3.835 0.68 3.835 1.25 5.845 1.25 5.845 0.68 6.075 0.68 6.075 1.25 8.085 1.25 8.085 0.68 8.315 0.68 8.315 1.25 9.32 1.25 9.32 2.27 11.05 2.27 11.05 2.5 9.32 2.5 9.32 4.09 4.72 4.09  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or4_4
