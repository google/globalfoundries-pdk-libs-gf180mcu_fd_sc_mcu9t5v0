# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 25.2 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.51 1.77 4.07 1.77 4.07 2.71 3.51 2.71  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.32 1.53 2.32 1.53 2.71 0.71 2.71  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER METAL1 ;
        POLYGON 18.63 1.21 18.89 1.21 18.89 2.265 19.11 2.265 19.11 2.605 18.63 2.605  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 2.32 2.65 2.32 2.65 2.71 1.83 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.865 2.32 7.69 2.32 7.69 2.71 6.865 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER METAL1 ;
        POLYGON 23.605 0.845 23.93 0.845 23.93 4.05 23.605 4.05  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.44 4.59 1.44 3.4 1.67 3.4 1.67 4.59 5.16 4.59 5.16 3.76 5.39 3.76 5.39 4.59 7.36 4.59 7.36 3.86 7.59 3.86 7.59 4.59 9.48 4.59 9.975 4.59 12.28 4.59 12.28 3.56 12.51 3.56 12.51 4.59 14.54 4.59 14.54 3.56 14.77 3.56 14.77 4.59 16.33 4.59 18.44 4.59 18.44 3.295 18.67 3.295 18.67 4.59 19.69 4.59 20.48 4.59 20.48 3.24 20.71 3.24 20.71 4.59 22.585 4.59 22.585 3.24 22.815 3.24 22.815 4.59 23.255 4.59 24.625 4.59 24.625 3.24 24.855 3.24 24.855 4.59 25.2 4.59 25.2 5.49 23.255 5.49 19.69 5.49 16.33 5.49 9.975 5.49 9.48 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 25.2 -0.45 25.2 0.45 24.955 0.45 24.955 1.165 24.725 1.165 24.725 0.45 22.715 0.45 22.715 1.165 22.485 1.165 22.485 0.45 20.61 0.45 20.61 1.48 20.38 1.48 20.38 0.45 12.51 0.45 12.51 1.22 12.28 1.22 12.28 0.45 7.59 0.45 7.59 1.17 7.36 1.17 7.36 0.45 5.775 0.45 5.775 0.575 5.545 0.575 5.545 0.45 1.67 0.45 1.67 1.48 1.44 1.48 1.44 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.42 2.94 2.88 2.94 2.88 2.09 0.32 2.09 0.32 1.14 0.55 1.14 0.55 1.86 3.11 1.86 3.11 2.94 4.4 2.94 4.4 2.84 4.68 2.84 4.68 2.265 4.91 2.265 4.91 3.07 4.59 3.07 4.59 3.17 0.65 3.17 0.65 4.05 0.42 4.05  ;
        POLYGON 6.34 2.875 6.57 2.875 6.57 2.94 7.92 2.94 7.92 2.09 6.24 2.09 6.24 1.26 6.47 1.26 6.47 1.86 8.15 1.86 8.15 3.17 6.57 3.17 6.57 3.215 6.34 3.215  ;
        POLYGON 3.4 0.805 6.14 0.805 6.14 0.8 6.93 0.8 6.93 1.4 7.82 1.4 7.82 0.68 9.43 0.68 9.43 1.22 9.2 1.22 9.2 0.91 8.05 0.91 8.05 1.63 6.7 1.63 6.7 1.03 6.19 1.03 6.19 1.035 3.63 1.035 3.63 1.48 3.4 1.48  ;
        POLYGON 3.4 3.4 4.78 3.4 4.78 3.3 5.82 3.3 5.82 3.445 7.08 3.445 7.08 3.4 8.05 3.4 8.05 3.915 9.25 3.915 9.25 3.09 9.48 3.09 9.48 4.145 7.82 4.145 7.82 3.63 7.22 3.63 7.22 3.675 5.605 3.675 5.605 3.53 4.97 3.53 4.97 3.63 3.63 3.63 3.63 4.21 3.4 4.21  ;
        POLYGON 8.38 1.14 8.71 1.14 8.71 2.32 9.975 2.32 9.975 2.55 8.61 2.55 8.61 3.685 8.38 3.685  ;
        POLYGON 10.32 1.11 10.55 1.11 10.55 2.085 11.555 2.085 11.555 2.055 13.225 2.055 13.225 2.285 11.67 2.285 11.67 2.315 10.55 2.315 10.55 3.73 10.32 3.73  ;
        POLYGON 10.845 1.595 12.74 1.595 12.74 0.68 15.265 0.68 15.265 0.91 12.97 0.91 12.97 1.825 11.185 1.825 11.185 1.855 10.845 1.855  ;
        POLYGON 11.785 2.515 14.54 2.515 14.54 1.14 14.77 1.14 14.77 2.515 15.89 2.515 15.89 3.685 15.66 3.685 15.66 2.745 13.75 2.745 13.75 3.73 13.52 3.73 13.52 2.745 11.785 2.745  ;
        POLYGON 10.9 3.1 12.97 3.1 12.97 3.96 14.08 3.96 14.08 3.1 15.43 3.1 15.43 3.975 16.33 3.975 16.33 4.315 15.2 4.315 15.2 3.33 14.31 3.33 14.31 4.19 12.74 4.19 12.74 3.33 11.13 3.33 11.13 4.36 10.9 4.36  ;
        POLYGON 17.72 2.835 18.17 2.835 18.17 1.655 16.78 1.655 16.78 1.315 18.4 1.315 18.4 2.835 19.69 2.835 19.69 4.05 19.46 4.05 19.46 3.065 17.95 3.065 17.95 3.845 17.72 3.845  ;
        POLYGON 15.66 1.14 16.32 1.14 16.32 0.75 19.35 0.75 19.35 1.71 20.73 1.71 20.73 2.32 21.385 2.32 21.385 2.55 20.5 2.55 20.5 1.94 19.12 1.94 19.12 0.98 16.55 0.98 16.55 1.885 16.91 1.885 16.91 3.845 16.68 3.845 16.68 2.115 16.32 2.115 16.32 1.48 15.66 1.48  ;
        POLYGON 20.04 2.265 20.27 2.265 20.27 2.78 21.68 2.78 21.68 0.845 21.91 0.845 21.91 2.78 23.025 2.78 23.025 2.265 23.255 2.265 23.255 3.01 21.91 3.01 21.91 4.05 21.68 4.05 21.68 3.01 20.04 3.01  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2
