# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.16 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.755 5.805 1.755 5.805 2.17 6.64 2.17 6.64 2.4 5.575 2.4 5.575 1.985 4.89 1.985 4.89 2.15 3.85 2.15 3.85 2.4 3.51 2.4  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.545 2.215 1.775 2.215 1.775 2.63 5.115 2.63 5.115 2.215 5.345 2.215 5.345 2.63 6.87 2.63 6.87 2.215 8.725 2.215 8.725 2.86 1.545 2.86  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.86 2.27 10.2 2.27 10.2 2.73 13.505 2.73 13.505 2.215 13.735 2.215 13.735 2.73 18.96 2.73 18.96 2.27 19.45 2.27 19.45 2.96 9.86 2.96  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.52 1.755 14.42 1.755 14.42 2.27 16.5 2.27 16.5 2.5 14.19 2.5 14.19 2.15 13.96 2.15 13.96 1.985 12.86 1.985 12.86 2.5 12.52 2.5  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.682 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.085 1.31 2.955 1.31 2.955 0.68 3.185 0.68 3.185 1.18 18.67 1.18 18.67 1.525 3.04 1.525 3.04 1.54 1.315 1.54 1.315 3.09 8.285 3.09 8.285 3.9 8.055 3.9 8.055 3.32 6.245 3.32 6.245 3.9 5.75 3.9 5.75 3.32 4.205 3.32 4.205 3.9 3.975 3.9 3.975 3.32 2.165 3.32 2.165 3.9 1.935 3.9 1.935 3.32 1.085 3.32  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 11.475 4.59 11.475 3.65 11.705 3.65 11.705 4.59 16.795 4.59 16.795 3.65 17.025 3.65 17.025 4.59 19.685 4.59 20.16 4.59 20.16 5.49 19.685 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 20.16 -0.45 20.16 0.45 19.735 0.45 19.735 1.035 19.505 1.035 19.505 0.45 17.34 0.45 17.34 0.95 17 0.95 17 0.45 14.68 0.45 14.68 0.95 14.34 0.95 14.34 0.45 12.02 0.45 12.02 0.95 11.68 0.95 11.68 0.45 9.36 0.45 9.36 0.95 9.02 0.95 9.02 0.45 5.225 0.45 5.225 0.695 4.995 0.695 4.995 0.45 0.905 0.45 0.905 1.165 0.675 1.165 0.675 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.915 3.55 1.145 3.55 1.145 4.13 2.955 4.13 2.955 3.55 3.185 3.55 3.185 4.13 4.995 4.13 4.995 3.55 5.225 3.55 5.225 4.13 7.035 4.13 7.035 3.55 7.265 3.55 7.265 4.13 9.075 4.13 9.075 3.19 19.685 3.19 19.685 4.36 19.455 4.36 19.455 3.42 14.365 3.42 14.365 4.36 14.135 4.36 14.135 3.42 9.305 3.42 9.305 4.36 0.915 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_4
