# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.79 2.33 3.29 2.33 4.36 2.33 4.36 2.71 3.29 2.71 1.79 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.77 2.33 1.11 2.33 1.11 2.94 3.29 2.94 4.63 2.94 4.63 2.33 5.43 2.33 5.43 2.71 4.86 2.71 4.86 3.17 3.29 3.17 0.77 3.17  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 3.45 7.665 3.45 7.665 0.845 7.895 0.845 7.895 1.885 9.905 1.885 9.905 0.845 10.135 0.845 10.135 4.36 9.855 4.36 9.855 2.115 7.895 2.115 7.895 4.36 7.43 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.86 0.475 3.86 0.475 4.59 2.285 4.59 2.285 3.86 2.515 3.86 2.515 4.59 3.29 4.59 5.725 4.59 5.725 3.86 5.955 3.86 5.955 4.59 6.645 4.59 6.645 3.86 6.875 3.86 6.875 4.59 7.315 4.59 8.735 4.59 8.735 3.86 8.965 3.86 8.965 4.59 10.925 4.59 10.925 3.86 11.155 3.86 11.155 4.59 11.76 4.59 11.76 5.49 7.315 5.49 3.29 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 11.255 0.45 11.255 1.655 11.025 1.655 11.025 0.45 9.015 0.45 9.015 1.655 8.785 1.655 8.785 0.45 6.775 0.45 6.775 1.165 6.545 1.165 6.545 0.45 2.57 0.45 2.57 1.595 2.23 1.595 2.23 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 1.365 0.53 1.365 0.53 1.87 3.29 1.87 3.29 2.1 0.42 2.1 0.42 3.4 1.495 3.4 1.495 4.065 1.265 4.065 1.265 3.63 0.19 3.63  ;
        POLYGON 3.585 0.83 6.055 0.83 6.055 1.64 5.825 1.64 5.825 1.06 3.815 1.06 3.815 1.65 3.585 1.65  ;
        POLYGON 3.635 3.4 5.66 3.4 5.66 2.1 4.705 2.1 4.705 1.31 4.935 1.31 4.935 1.87 7.315 1.87 7.315 2.21 5.89 2.21 5.89 3.63 3.865 3.63 3.865 4.36 3.635 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_4
