# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 1.77 5.45 1.77 5.45 2.15 4.63 2.15  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 1.77 2.65 1.77 2.65 2.71 2.39 2.71  ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.225 1.38 3.455 1.38 3.455 2.475 5.75 2.475 5.75 1.77 6.035 1.77 6.035 3.27 5.75 3.27 5.75 2.705 3.225 2.705  ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 0.72 0.575 0.72 0.575 4.235 0.15 4.235  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 2.97 1.595 2.97 1.595 4.59 3.835 4.59 5.31 4.59 5.31 3.48 5.65 3.48 5.65 4.59 6.815 4.59 7.28 4.59 7.28 5.49 6.815 5.49 3.835 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 5.695 0.45 5.695 0.99 5.465 0.99 5.465 0.45 1.595 0.45 1.595 1.06 1.365 1.06 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.16 3.545 3.605 3.545 3.605 2.965 3.835 2.965 3.835 3.775 1.93 3.775 1.93 2.055 0.87 2.055 0.87 1.825 1.93 1.825 1.93 0.775 3.79 0.775 3.79 1.005 2.16 1.005  ;
        POLYGON 3.945 1.31 6.585 1.31 6.585 0.72 6.815 0.72 6.815 3.775 6.385 3.775 6.385 1.54 4.175 1.54 4.175 2.11 3.945 2.11  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_1
