* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I B1:I B2:I C:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(((A1 * A2) + (B1 * B2)) + C)
M_i_2_1 VSS C ZN VPW nfet_05v0 W=0.790000U L=0.600000U
M_i_4_1 net_1_0 B2 VSS VPW nfet_05v0 W=1.185000U L=0.600000U
M_i_3_1 ZN B1 net_1_0 VPW nfet_05v0 W=1.185000U L=0.600000U
M_i_3_0 net_1_1 B1 ZN VPW nfet_05v0 W=1.185000U L=0.600000U
M_i_4_0 VSS B2 net_1_1 VPW nfet_05v0 W=1.185000U L=0.600000U
M_i_2_0 ZN C VSS VPW nfet_05v0 W=0.790000U L=0.600000U
M_i_0_1 net_0_0 A1 ZN VPW nfet_05v0 W=1.185000U L=0.600000U
M_i_1_1 VSS A2 net_0_0 VPW nfet_05v0 W=1.185000U L=0.600000U
M_i_1_0 net_0_1 A2 VSS VPW nfet_05v0 W=1.185000U L=0.600000U
M_i_0_0 ZN A1 net_0_1 VPW nfet_05v0 W=1.185000U L=0.600000U
M_i_7_1 net_3 C net_2 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_1 VDD B2 net_3 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8_1 net_3 B1 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8_0 VDD B1 net_3 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_0 net_3 B2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_7_0 net_2 C net_3 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_5_1 ZN A1 net_2 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_1 net_2 A2 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_0 ZN A2 net_2 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_5_0 net_2 A1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
