# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.63 2.27 5.5 2.27 5.5 2.71 4.63 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.51 1.77 3.77 1.77 3.77 1.81 6.275 1.81 6.275 2.215 7.685 2.215 7.685 2.555 6.045 2.555 6.045 2.04 4.38 2.04 4.38 2.5 4.04 2.5 4.04 2.15 3.51 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.055 2.215 3.285 2.215 3.285 2.94 7.99 2.94 7.99 2.215 8.755 2.215 8.755 2.71 8.22 2.71 8.22 3.17 3.055 3.17  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.675 2.215 0.97 2.215 0.97 2.71 0.675 2.71  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.13145 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.365 3.4 8.985 3.4 8.985 1.935 6.505 1.935 6.505 1.58 3.935 1.58 3.935 1.54 3.605 1.54 3.605 1.14 4.065 1.14 4.065 1.35 5.845 1.35 5.845 1.14 6.735 1.14 6.735 1.705 7.43 1.705 7.43 1.14 8.315 1.14 8.315 1.705 9.215 1.705 9.215 3.63 6.025 3.63 6.025 4.36 5.795 4.36 5.795 3.63 1.595 3.63 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.86 0.525 3.86 0.525 4.59 2.385 4.59 2.385 3.86 2.615 3.86 2.615 4.59 9.105 4.59 9.105 3.86 9.335 3.86 9.335 4.59 9.67 4.59 10.08 4.59 10.08 5.49 9.67 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 1.595 0.45 1.595 1.525 1.365 1.525 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 1.755 2.485 1.755 2.485 0.68 9.67 0.68 9.67 1.655 9.44 1.655 9.44 0.91 7.195 0.91 7.195 1.185 6.965 1.185 6.965 0.91 4.955 0.91 4.955 1.12 4.725 1.12 4.725 0.91 2.715 0.91 2.715 1.985 0.245 1.985  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_2
