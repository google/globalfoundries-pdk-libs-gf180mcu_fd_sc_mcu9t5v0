# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__and4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 13.44 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.79 1.77 3.89 1.77 3.89 2.15 2.79 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.825 2.38 4.52 2.38 4.52 1.77 6.03 1.77 6.03 2.15 4.75 2.15 4.75 2.61 2.825 2.61  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.975 1.21 2.09 1.21 2.09 1.31 6.49 1.31 6.49 1.83 7.105 1.83 7.105 2.06 6.26 2.06 6.26 1.54 2.145 1.54 2.145 2.06 0.975 2.06  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.33 0.97 2.33 0.97 2.84 4.98 2.84 4.98 2.47 8.125 2.47 8.125 2.7 5.21 2.7 5.21 3.07 0.115 3.07  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.54 2.92 10.55 2.92 11.77 2.92 11.77 1.6 9.485 1.6 9.485 0.9 12.21 0.9 12.21 3.64 10.55 3.64 9.54 3.64  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.26 4.59 0.26 3.325 0.49 3.325 0.49 4.59 2.3 4.59 2.3 3.795 2.53 3.795 2.53 4.59 4.34 4.59 4.34 3.795 4.57 3.795 4.57 4.59 6.38 4.59 6.38 3.795 6.61 3.795 6.61 4.59 8.42 4.59 8.42 3.795 8.65 3.795 8.65 4.59 10.55 4.59 10.64 4.59 10.64 3.875 10.87 3.875 10.87 4.59 12.68 4.59 12.68 3.875 12.91 3.875 12.91 4.59 13.44 4.59 13.44 5.49 10.55 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 13.44 -0.45 13.44 0.45 13.13 0.45 13.13 1.165 12.9 1.165 12.9 0.45 10.945 0.45 10.945 0.64 10.605 0.64 10.605 0.45 8.65 0.45 8.65 0.695 8.42 0.695 8.42 0.45 0.49 0.45 0.49 1.165 0.26 1.165 0.26 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.28 3.3 5.4 3.3 5.4 3.2 8.86 3.2 8.86 1.26 6.715 1.26 6.715 1.08 4.285 1.08 4.285 0.85 6.94 0.85 6.94 1.03 9.09 1.03 9.09 1.975 10.55 1.975 10.55 2.315 9.09 2.315 9.09 3.43 7.63 3.43 7.63 4.01 7.4 4.01 7.4 3.43 5.59 3.43 5.59 4.11 5.36 4.11 5.36 3.53 3.55 3.53 3.55 4.11 3.32 4.11 3.32 3.53 1.51 3.53 1.51 4.11 1.28 4.11  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_4
