# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__and2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.806 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.15 0.97 2.15 0.97 2.96 0.71 2.96 0.71 2.71 0.115 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.806 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.15 2.715 2.15 2.715 2.71 2.06 2.71 2.06 2.96 1.83 2.96  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 0.845 3.855 0.845 3.855 3.685 3.51 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 4.345 0.475 4.345 0.475 4.59 2.285 4.59 2.285 4.345 2.515 4.345 2.515 4.59 3.175 4.59 4.48 4.59 4.48 5.49 3.175 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 2.735 0.45 2.735 1.165 2.505 1.165 2.505 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.21 3.885 2.945 3.885 2.945 1.625 0.19 1.625 0.19 1.37 0.53 1.37 0.53 1.395 3.175 1.395 3.175 4.115 1.55 4.115 1.55 4.17 1.21 4.17  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and2_1
