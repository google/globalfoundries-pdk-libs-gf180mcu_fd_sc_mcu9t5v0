# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi22_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.96 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.75 1.72 7.21 1.72 7.21 2.315 5.75 2.315  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.95 1.83 5.51 1.83 5.51 2.56 7.86 2.56 7.86 2.18 8.27 2.18 8.27 2.79 4.95 2.79  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.22 1.21 2.09 1.21 2.09 2.06 1.65 2.06 1.65 1.63 1.22 1.63  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.69 1.77 0.97 1.77 0.97 2.29 4.03 2.29 4.03 2.52 0.69 2.52  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.3222 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.72 3.02 7.615 3.02 7.615 3.83 7.385 3.83 7.385 3.25 5.575 3.25 5.575 3.83 4.345 3.83 4.345 1.49 4.34 1.49 4.34 1.105 2.55 1.105 2.55 1.49 2.32 1.49 2.32 0.68 2.55 0.68 2.55 0.875 6.365 0.875 6.365 0.68 6.595 0.68 6.595 1.49 6.365 1.49 6.365 1.105 4.72 1.105  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.875 1.495 3.875 1.495 4.59 3.305 4.59 3.305 3.875 3.535 3.875 3.535 4.59 8.635 4.59 8.96 4.59 8.96 5.49 8.635 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 8.96 -0.45 8.96 0.45 8.635 0.45 8.635 1.165 8.405 1.165 8.405 0.45 4.61 0.45 4.61 0.64 4.27 0.64 4.27 0.45 0.475 0.45 0.475 1.165 0.245 1.165 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 3.415 4.025 3.415 4.025 4.06 6.365 4.06 6.365 3.48 6.595 3.48 6.595 4.06 8.405 4.06 8.405 3.48 8.635 3.48 8.635 4.29 3.795 4.29 3.795 3.645 2.515 3.645 2.515 4.225 2.285 4.225 2.285 3.645 0.475 3.645 0.475 4.225 0.245 4.225  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi22_2
