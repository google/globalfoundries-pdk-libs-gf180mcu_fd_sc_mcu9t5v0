# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.68 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.165 1.72 4.33 1.72 4.33 2.18 4.575 2.18 4.575 2.52 4.07 2.52 4.07 1.95 2.395 1.95 2.395 2.52 2.165 2.52  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.025 2.18 1.255 2.18 1.255 3.21 3.555 3.21 5.19 3.21 5.19 2.18 5.595 2.18 5.595 3.44 3.555 3.44 1.025 3.44  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.31 2.77 9.86 2.77 10.23 2.77 10.23 2.31 10.93 2.31 10.93 2.54 10.49 2.54 10.49 3 9.86 3 8.31 3  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.772 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.015 3.155 13.685 3.155 13.915 3.155 13.915 1.945 12.965 1.945 12.965 0.845 13.29 0.845 13.29 1.715 15.205 1.715 15.205 0.845 15.435 0.845 15.435 1.945 14.145 1.945 14.145 3.155 15.385 3.155 15.385 4.36 15.155 4.36 15.155 3.385 13.685 3.385 13.245 3.385 13.245 4.36 13.015 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.605 4.59 2.605 3.67 2.835 3.67 2.835 4.59 3.555 4.59 6.23 4.59 8.805 4.59 8.805 3.615 9.035 3.615 9.035 4.59 9.86 4.59 12.475 4.59 13.685 4.59 14.035 4.59 14.035 3.615 14.265 3.615 14.265 4.59 15.68 4.59 15.68 5.49 13.685 5.49 12.475 5.49 9.86 5.49 6.23 5.49 3.555 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 15.68 -0.45 15.68 0.45 14.315 0.45 14.315 1.485 14.085 1.485 14.085 0.45 12.475 0.45 12.475 1.16 12.245 1.16 12.245 0.45 9.315 0.45 9.315 1.18 9.085 1.18 9.085 0.45 6.895 0.45 6.895 1.185 6.665 1.185 6.665 0.45 6.175 0.45 6.175 1.185 5.945 1.185 5.945 0.45 2.835 0.45 2.835 1.185 2.605 1.185 2.605 0.45 0.595 0.45 0.595 1.185 0.365 1.185 0.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.465 1.72 1.485 1.72 1.485 0.845 1.715 0.845 1.715 2.75 3.325 2.75 3.325 2.18 3.555 2.18 3.555 2.98 1.485 2.98 1.485 1.95 0.695 1.95 0.695 3.955 0.465 3.955  ;
        POLYGON 3.905 3.67 4.135 3.67 4.135 4.13 6.23 4.13 6.23 4.36 3.905 4.36  ;
        POLYGON 6.765 2.75 7.785 2.75 7.785 1.145 8.015 1.145 8.015 2.31 9.86 2.31 9.86 2.54 8.015 2.54 8.015 2.98 6.995 2.98 6.995 4.36 6.765 4.36  ;
        POLYGON 4.87 3.67 5.825 3.67 5.825 2.29 7.205 2.29 7.205 1.645 4.55 1.645 4.55 1.13 3.85 1.13 3.85 0.9 4.78 0.9 4.78 1.415 7.205 1.415 7.205 0.685 8.475 0.685 8.475 1.85 11.895 1.85 11.895 2.52 11.665 2.52 11.665 2.08 8.245 2.08 8.245 0.915 7.435 0.915 7.435 2.52 6.055 2.52 6.055 3.9 4.87 3.9  ;
        POLYGON 10.15 3.55 12.475 3.55 12.475 4.36 12.245 4.36 12.245 3.9 10.15 3.9  ;
        POLYGON 11.17 2.93 12.125 2.93 12.125 1.62 10.205 1.62 10.205 0.845 10.435 0.845 10.435 1.39 12.355 1.39 12.355 2.18 13.685 2.18 13.685 2.52 12.355 2.52 12.355 3.16 11.17 3.16  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_2
