# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.64 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.87 2.33 2.09 2.33 2.09 2.71 0.87 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.547 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.75 1.75 6.115 1.75 6.115 2.15 5.75 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.9952 ;
    PORT
      LAYER METAL1 ;
        POLYGON 7.895 2.91 9.045 2.91 9.045 1.65 7.865 1.65 7.865 0.84 8.095 0.84 8.095 1.39 10.105 1.39 10.105 0.84 10.335 0.84 10.335 1.65 9.39 1.65 9.39 2.91 10.165 2.91 10.165 3.72 9.935 3.72 9.935 3.14 8.125 3.14 8.125 3.72 7.895 3.72  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.845 1.595 3.845 1.595 4.59 4.655 4.59 4.655 4.035 4.885 4.035 4.885 4.59 6.695 4.59 6.695 3.565 6.925 3.565 6.925 4.59 7.665 4.59 8.915 4.59 8.915 3.88 9.145 3.88 9.145 4.59 10.64 4.59 10.64 5.49 7.665 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 10.64 -0.45 10.64 0.45 9.215 0.45 9.215 1.16 8.985 1.16 8.985 0.45 6.85 0.45 6.85 0.68 6.51 0.68 6.51 0.45 4.61 0.45 4.61 0.68 4.27 0.68 4.27 0.45 1.595 0.45 1.595 1.165 1.365 1.165 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.845 0.475 0.845 0.475 1.83 2.55 1.83 2.55 2.47 3.65 2.47 3.65 2.7 2.32 2.7 2.32 2.06 0.575 2.06 0.575 3.685 0.245 3.685  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.91 6.575 0.91 6.575 1.825 7.665 1.825 7.665 2.055 6.345 2.055 6.345 1.14 3.32 1.14 3.32 1.83 4.165 1.83 4.165 3.215 3.935 3.215 3.935 2.06 3.09 2.06 3.09 1.49 2.485 1.49  ;
        POLYGON 2.915 2.93 3.145 2.93 3.145 3.51 5.675 3.51 5.675 2.695 5.29 2.695 5.29 1.6 3.55 1.6 3.55 1.37 5.52 1.37 5.52 2.465 7.665 2.465 7.665 2.695 5.905 2.695 5.905 3.74 2.915 3.74  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_3
