# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi221_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.225 2.47 10.165 2.47 10.165 1.21 10.49 1.21 10.49 2.7 7.225 2.7  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.3 1.21 8.47 1.21 8.47 2.115 8.24 2.115 8.24 1.59 7.3 1.59  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 1.665 3.845 1.665 3.845 2.18 2.945 2.18  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.89 2.44 4.49 2.44 4.49 2.205 5.48 2.205 5.48 2.67 1.89 2.67  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.715 1.915 2.485 1.915 2.485 1.205 4.89 1.205 4.89 1.52 6.37 1.52 6.37 1.75 4.63 1.75 4.63 1.435 2.715 1.435 2.715 2.145 1.01 2.145 1.01 2.785 0.715 2.785  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.11125 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.245 1.315 0.475 1.315 0.475 1.455 2.025 1.455 2.025 0.745 5.35 0.745 5.35 1.06 6.765 1.06 6.765 0.92 6.995 0.92 6.995 3.02 10.88 3.02 10.88 0.845 11.11 0.845 11.11 3.83 9.76 3.83 9.76 3.25 7.95 3.25 7.95 3.83 7.72 3.83 7.72 3.25 6.765 3.25 6.765 1.29 5.12 1.29 5.12 0.975 2.255 0.975 2.255 1.685 0.245 1.685  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.33 4.59 2.33 4.4 2.67 4.4 2.67 4.59 4.39 4.59 4.39 4.4 4.73 4.4 4.73 4.59 11.065 4.59 11.76 4.59 11.76 5.49 11.065 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 9.15 0.45 9.15 1.3 8.92 1.3 8.92 0.45 5.81 0.45 5.81 0.83 5.58 0.83 5.58 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.9 1.595 2.9 1.595 3.48 3.405 3.48 3.405 2.9 3.635 2.9 3.635 3.48 5.465 3.48 5.465 2.9 5.695 2.9 5.695 3.71 1.365 3.71  ;
        POLYGON 0.345 3.36 0.575 3.36 0.575 3.94 6.665 3.94 6.665 3.48 6.895 3.48 6.895 4.06 8.74 4.06 8.74 3.48 8.97 3.48 8.97 4.06 11.065 4.06 11.065 4.29 6.665 4.29 6.665 4.17 0.345 4.17  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi221_2
