# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__and3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.125 2.74 1.145 2.74 1.145 3.345 0.125 3.345  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.82 2.74 2.725 2.74 2.725 3.375 1.82 3.375  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.761 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.565 1.77 2.955 1.77 2.955 2.15 0.565 2.15  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.63 0.845 4.995 0.845 4.995 3.83 4.63 3.83  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 4.345 1.495 4.345 1.495 4.59 3.645 4.59 3.645 4.345 3.875 4.345 3.875 4.59 4.315 4.59 5.6 4.59 5.6 5.49 4.315 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 3.875 0.45 3.875 1.35 3.645 1.35 3.645 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 3.885 3.185 3.885 3.185 0.98 0.475 0.98 0.475 1.355 0.245 1.355 0.245 0.75 3.415 0.75 3.415 1.775 4.315 1.775 4.315 2.115 3.415 2.115 3.415 4.315 2.285 4.315 2.285 4.115 0.475 4.115 0.475 4.315 0.245 4.315  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and3_1
