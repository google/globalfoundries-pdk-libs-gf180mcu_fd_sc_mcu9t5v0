# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.72 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.965 2.315 4.01 2.315 4.01 2.545 3.77 2.545 3.77 2.71 2.965 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER METAL1 ;
        POLYGON 16.3 2.33 17.21 2.33 17.21 2.89 16.3 2.89  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.71 2.89 14.825 2.89 14.825 2.47 15.055 2.47 15.055 3.27 14.71 3.27  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.48 1.58 2.48 1.58 3.27 0.71 3.27  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 19.125 0.845 19.45 0.845 19.45 3.685 19.125 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.96 1.495 3.96 1.495 4.59 2.055 4.59 3.005 4.59 3.005 3.56 3.235 3.56 3.235 4.59 4.835 4.59 7.245 4.59 7.245 4.49 7.475 4.49 7.475 4.59 10.445 4.59 10.445 4.49 10.675 4.49 10.675 4.59 12.49 4.59 14.33 4.59 14.33 4.005 14.67 4.005 14.67 4.59 16.37 4.59 16.37 4.005 16.71 4.005 16.71 4.59 18.135 4.59 18.465 4.59 18.465 3.48 18.695 3.48 18.695 4.59 18.895 4.59 20.205 4.59 20.205 3.875 20.435 3.875 20.435 4.59 20.72 4.59 20.72 5.49 18.895 5.49 18.135 5.49 12.49 5.49 4.835 5.49 2.055 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 20.72 -0.45 20.72 0.45 20.475 0.45 20.475 1.165 20.245 1.165 20.245 0.45 16.59 0.45 16.59 1.225 16.36 1.225 16.36 0.45 8.815 0.45 8.815 1.425 8.585 1.425 8.585 0.45 3.515 0.45 3.515 1.425 3.285 1.425 3.285 0.45 1.615 0.45 1.615 1.225 1.385 1.225 1.385 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 3.39 0.475 3.39 0.475 3.5 1.825 3.5 1.825 1.74 0.265 1.74 0.265 1.315 0.495 1.315 0.495 1.51 2.055 1.51 2.055 3.73 0.245 3.73  ;
        POLYGON 4.025 2.775 4.405 2.775 4.405 1.315 4.635 1.315 4.635 3.005 4.255 3.005 4.255 3.73 4.025 3.73  ;
        POLYGON 2.285 1.315 2.735 1.315 2.735 3.1 3.695 3.1 3.695 4.02 4.835 4.02 4.835 4.36 3.465 4.36 3.465 3.33 2.515 3.33 2.515 3.75 2.285 3.75  ;
        POLYGON 6.065 3.35 8.715 3.35 8.715 3.8 6.065 3.8  ;
        POLYGON 5.045 2.685 5.525 2.685 5.525 1.315 5.755 1.315 5.755 2.685 9.265 2.685 9.265 2.575 9.495 2.575 9.495 2.915 5.275 2.915 5.275 3.73 5.045 3.73  ;
        POLYGON 9.955 3.57 11.625 3.57 11.625 2.875 11.855 2.875 11.855 3.8 9.205 3.8 9.205 3.46 9.725 3.46 9.725 2.345 7.035 2.345 7.035 2.455 6.805 2.455 6.805 2.115 10.545 2.115 10.545 1.315 10.775 1.315 10.775 2.345 9.955 2.345  ;
        POLYGON 5.57 4.03 12.49 4.03 12.49 4.26 5.91 4.26 5.91 4.305 5.57 4.305  ;
        POLYGON 5.985 1.655 10.085 1.655 10.085 0.68 13.525 0.68 13.525 2.275 13.295 2.275 13.295 0.91 10.315 0.91 10.315 1.885 6.215 1.885 6.215 2.115 5.985 2.115  ;
        POLYGON 12.785 1.315 13.015 1.315 13.015 2.505 14.265 2.505 14.265 1.315 14.63 1.315 14.63 2.01 15.635 2.01 15.635 3.27 15.405 3.27 15.405 2.24 14.495 2.24 14.495 2.735 13.895 2.735 13.895 3.215 13.665 3.215 13.665 2.735 12.785 2.735  ;
        POLYGON 11.665 1.315 11.895 1.315 11.895 2.415 12.315 2.415 12.315 2.965 12.875 2.965 12.875 3.545 17.905 3.545 17.905 2.47 18.135 2.47 18.135 3.775 12.645 3.775 12.645 3.195 12.085 3.195 12.085 2.645 11.665 2.645  ;
        POLYGON 15.865 1.83 18.32 1.83 18.32 1.315 18.55 1.315 18.55 1.975 18.895 1.975 18.895 2.315 18.32 2.315 18.32 2.06 17.675 2.06 17.675 3.27 17.445 3.27 17.445 2.06 15.865 2.06  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1
