* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I A3:I B:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(((A1 + A2) + A3) * B)
M_i_3 net_0 B VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1 net_0 A2 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 ZN A3 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_7 ZN B VDD VNW pmos_5p0 W=1.645000U L=0.500000U
M_i_4 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 net_2 A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 VDD A3 net_2 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
