# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 29.12 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.51 1.77 3.77 1.77 3.77 2.71 3.51 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123 ;
    PORT
      LAYER METAL1 ;
        POLYGON 21.43 2.215 21.69 2.215 21.69 3.27 21.43 3.27  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 2.27 0.97 2.27 0.97 2.71 0.15 2.71  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER METAL1 ;
        POLYGON 19.13 2.95 19.655 2.95 19.655 2.74 20.01 2.74 20.01 3.27 19.13 3.27  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.27 2.27 2.09 2.27 2.09 2.71 1.27 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.75 2.89 6.28 2.89 6.28 2.53 6.57 2.53 6.57 3.27 5.75 3.27  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER METAL1 ;
        POLYGON 24.85 2.89 25.25 2.89 25.25 0.845 25.48 0.845 25.48 2.89 27.49 2.89 27.49 0.845 27.72 0.845 27.72 3.12 26.73 3.12 26.73 3.44 27.12 3.44 27.12 4.25 26.47 4.25 26.47 3.12 25.08 3.12 25.08 4.25 24.85 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.44 1.495 3.44 1.495 4.59 4.95 4.59 4.95 4.56 5.29 4.56 5.29 4.59 6.885 4.59 6.885 4.56 7.225 4.56 7.225 4.59 9.13 4.59 9.57 4.59 9.61 4.59 12.12 4.59 12.12 4.51 12.35 4.51 12.35 4.59 15.32 4.59 15.32 4.51 15.55 4.51 15.55 4.59 17.355 4.59 19.39 4.59 19.39 3.985 19.62 3.985 19.62 4.59 21.595 4.59 21.595 4.375 21.935 4.375 21.935 4.59 23.36 4.59 23.71 4.59 23.71 3.44 23.94 3.44 23.94 4.59 24.8 4.59 25.87 4.59 25.87 3.44 26.1 3.44 26.1 4.59 27.91 4.59 27.91 3.44 28.14 3.44 28.14 4.59 29.12 4.59 29.12 5.49 24.8 5.49 23.36 5.49 17.355 5.49 9.61 5.49 9.57 5.49 9.13 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 29.12 -0.45 29.12 0.45 28.84 0.45 28.84 1.65 28.61 1.65 28.61 0.45 26.6 0.45 26.6 1.65 26.37 1.65 26.37 0.45 24.36 0.45 24.36 1.525 24.13 1.525 24.13 0.45 21.22 0.45 21.22 1.255 20.99 1.255 20.99 0.45 13.69 0.45 13.69 1.535 13.46 1.535 13.46 0.45 7.69 0.45 7.69 1.38 7.46 1.38 7.46 0.45 5.675 0.45 5.675 0.53 5.445 0.53 5.445 0.45 1.595 0.45 1.595 1.535 1.365 1.535 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 2.94 2.445 2.94 2.445 2.04 0.245 2.04 0.245 1.195 0.475 1.195 0.475 1.81 2.675 1.81 2.675 2.94 4.605 2.94 4.605 2.215 4.835 2.215 4.835 3.17 0.475 3.17 0.475 4.25 0.245 4.25  ;
        POLYGON 5.7 3.5 7.6 3.5 7.6 2.3 6.34 2.3 6.34 1.22 6.57 1.22 6.57 2.07 7.83 2.07 7.83 3.84 5.7 3.84  ;
        POLYGON 3.025 3.44 3.255 3.44 3.255 4.1 8.9 4.1 8.9 3.065 9.13 3.065 9.13 4.33 3.025 4.33  ;
        POLYGON 8.18 2.325 8.58 2.325 8.58 1.22 8.81 1.22 8.81 2.215 9.57 2.215 9.57 2.555 8.41 2.555 8.41 3.87 8.18 3.87  ;
        POLYGON 3.325 0.76 7.03 0.76 7.03 1.61 8.12 1.61 8.12 0.76 9.61 0.76 9.61 1.535 9.38 1.535 9.38 0.99 8.35 0.99 8.35 1.84 6.8 1.84 6.8 0.99 3.555 0.99 3.555 1.535 3.325 1.535  ;
        POLYGON 10.94 3.44 13.59 3.44 13.59 3.78 10.94 3.78  ;
        POLYGON 9.92 2.985 10.5 2.985 10.5 1.195 10.73 1.195 10.73 2.98 14.75 2.98 14.75 3.32 14.52 3.32 14.52 3.21 10.55 3.21 10.55 3.215 10.15 3.215 10.15 3.875 9.92 3.875  ;
        POLYGON 14.08 3.44 14.31 3.44 14.31 3.55 15.64 3.55 15.64 2.565 11.92 2.565 11.92 2.225 15.64 2.225 15.64 1.195 15.87 1.195 15.87 3.44 16.86 3.44 16.86 3.78 14.08 3.78  ;
        POLYGON 10.445 4.05 17.355 4.05 17.355 4.28 10.445 4.28  ;
        POLYGON 11.08 1.765 15.18 1.765 15.18 0.68 18.68 0.68 18.68 2.22 18.34 2.22 18.34 0.91 15.41 0.91 15.41 1.995 11.31 1.995 11.31 2.115 11.08 2.115  ;
        POLYGON 17.88 1.195 18.11 1.195 18.11 2.45 19.03 2.45 19.03 1.145 19.26 1.145 19.26 2.28 20.64 2.28 20.64 3.685 20.41 3.685 20.41 2.51 19.255 2.51 19.255 2.68 18.9 2.68 18.9 3.295 18.67 3.295 18.67 2.68 17.88 2.68  ;
        POLYGON 16.76 1.195 16.99 1.195 16.99 2.945 17.88 2.945 17.88 3.525 20.08 3.525 20.08 3.915 23.13 3.915 23.13 2.215 23.36 2.215 23.36 4.145 19.85 4.145 19.85 3.755 17.65 3.755 17.65 3.175 16.76 3.175  ;
        POLYGON 20.795 1.755 23.41 1.755 23.41 0.845 23.64 0.845 23.64 1.755 24.8 1.755 24.8 2.555 24.57 2.555 24.57 1.985 22.9 1.985 22.9 3.685 22.67 3.685 22.67 1.985 21.135 1.985 21.135 2.11 20.795 2.11  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4
