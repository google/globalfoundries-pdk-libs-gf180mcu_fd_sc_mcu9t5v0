* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__dffnq_2 D CLKN Q VDD VNW VPW VSS
*.PININFO D:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G
M_tn9 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn16 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 VSS D net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn11 net2 cki net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn0 net5 ncki net11 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 VSS net10 net11 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn15 net10 net5 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn2 net0 ncki net10 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn3 net7 cki net0 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn4 VSS net1 net7 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn5 net1 net0 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6_7 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn6 Q net1 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp9 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp16 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp10 VDD D net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp11 net5 ncki net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp0 net4 cki net5 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp1 VDD net10 net4 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net10 net5 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net0 cki net10 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 net7 ncki net0 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 VDD net1 net7 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp3 net1 net0 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4_13 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4 Q net1 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
