* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__hold Z VDD VNW VPW VSS
*.PININFO Z:B VDD:P VNW:P VPW:P VSS:G
M_u7 VDD Z net8 VNW pmos_5p0 W=1.830000U L=0.500000U
M_u3 VSS Z net8 VPW nmos_5p0 W=1.320000U L=0.600000U
M_MU12 Z net8 VDD VNW pmos_5p0 W=0.360000U L=2.00000U
M_MU11 Z net8 VSS VPW nmos_5p0 W=0.360000U L=2.00000U
.ENDS
