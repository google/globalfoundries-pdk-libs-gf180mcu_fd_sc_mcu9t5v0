# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.6 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 1.77 3.895 1.77 3.895 2.15 2.945 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.38 1.675 14.41 1.675 14.41 2.15 13.38 2.15  ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.575 1.77 1.575 2.245 0.71 2.245  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.51 3.45 17.685 3.45 17.685 0.845 17.915 0.845 17.915 3.83 17.51 3.83  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.225 4.59 3.225 3.045 3.455 3.045 3.455 4.59 5.99 4.59 7.305 4.59 7.305 3.515 7.535 3.515 7.535 4.59 8.555 4.59 9.045 4.59 9.045 3.44 9.275 3.44 9.275 4.59 9.77 4.59 10.295 4.59 13.525 4.59 13.525 4.345 13.755 4.345 13.755 4.59 15.495 4.59 15.845 4.59 15.845 3.875 16.075 3.875 16.075 4.59 16.665 4.59 16.665 3.875 16.895 3.875 16.895 4.59 17.39 4.59 18.705 4.59 18.705 3.875 18.935 3.875 18.935 4.59 19.6 4.59 19.6 5.49 17.39 5.49 15.495 5.49 10.295 5.49 9.77 5.49 8.555 5.49 5.99 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.6 -0.45 19.6 0.45 19.035 0.45 19.035 1.165 18.805 1.165 18.805 0.45 16.795 0.45 16.795 1.165 16.565 1.165 16.565 0.45 13.655 0.45 13.655 1.31 13.425 1.31 13.425 0.45 8.655 0.45 8.655 1.31 8.425 1.31 8.425 0.45 3.435 0.45 3.435 1.31 3.205 1.31 3.205 0.45 1.65 0.45 1.65 1.08 1.31 1.08 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.875 1.805 2.875 1.805 1.54 0.245 1.54 0.245 1.19 0.475 1.19 0.475 1.31 2.035 1.31 2.035 3.105 0.575 3.105 0.575 3.685 0.345 3.685  ;
        POLYGON 4.245 1.31 4.555 1.31 4.555 3.685 4.245 3.685  ;
        POLYGON 2.385 1.19 2.715 1.19 2.715 2.585 3.915 2.585 3.915 4.03 5.99 4.03 5.99 4.26 3.685 4.26 3.685 2.815 2.615 2.815 2.615 3.685 2.385 3.685  ;
        POLYGON 6.285 2.92 8.555 2.92 8.555 3.73 8.325 3.73 8.325 3.15 6.515 3.15 6.515 3.73 6.285 3.73  ;
        POLYGON 5.265 1.31 5.675 1.31 5.675 2.46 9.77 2.46 9.77 2.69 5.495 2.69 5.495 3.685 5.265 3.685  ;
        POLYGON 6.81 2 10.065 2 10.065 1.31 10.295 1.31 10.295 4.08 10.065 4.08 10.065 2.23 6.81 2.23  ;
        POLYGON 6.07 1.825 6.35 1.825 6.35 1.54 9.605 1.54 9.605 0.85 11.875 0.85 11.875 3.15 11.645 3.15 11.645 1.08 10.755 1.08 10.755 2.11 10.525 2.11 10.525 1.08 9.835 1.08 9.835 1.77 6.58 1.77 6.58 2.055 6.07 2.055  ;
        POLYGON 12.285 1.31 12.535 1.31 12.535 3.61 12.285 3.61  ;
        POLYGON 11.185 1.31 11.415 1.31 11.415 3.27 11.42 3.27 11.42 3.85 15.265 3.85 15.265 2.415 15.495 2.415 15.495 4.08 11.185 4.08  ;
        POLYGON 12.81 2.38 14.805 2.38 14.805 1.955 15.845 1.955 15.845 0.845 16.075 0.845 16.075 1.83 17.39 1.83 17.39 2.185 15.035 2.185 15.035 2.61 14.775 2.61 14.775 3.215 14.545 3.215 14.545 2.61 12.81 2.61  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2
