# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai33_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai33_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 28.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.325 2.19 17.85 2.19 17.85 2.71 15.325 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.12 2.27 19.46 2.27 19.46 2.495 21.99 2.495 21.99 2.27 22.82 2.27 22.82 2.495 26.965 2.495 26.965 2.215 27.195 2.215 27.195 2.725 19.12 2.725  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.69 1.81 25.06 1.81 25.06 2.265 24.72 2.265 24.72 2.04 20.58 2.04 20.58 2.265 19.69 2.265  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.325 2.19 12.795 2.19 12.795 2.71 10.325 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.82 2.19 1.16 2.19 1.16 2.65 4.04 2.65 4.04 2.27 4.38 2.27 4.38 2.65 6.8 2.65 6.8 2.27 8.86 2.27 8.86 2.5 7.03 2.5 7.03 2.88 0.82 2.88  ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 4.84 1.77 4.84 2.19 6.57 2.19 6.57 2.42 4.61 2.42 4.61 2 2.17 2 2.17 2.42 1.83 2.42  ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.3823 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.325 2.955 27.425 2.955 27.425 1.53 15.27 1.53 15.27 1.3 17.51 1.3 17.51 1.14 17.85 1.14 17.85 1.3 19.75 1.3 19.75 1.14 20.09 1.14 20.09 1.3 21.99 1.3 21.99 1.14 22.33 1.14 22.33 1.3 24.23 1.3 24.23 1.14 24.57 1.14 24.57 1.3 27.655 1.3 27.655 3.185 17.745 3.185 17.745 3.46 17.515 3.46 17.515 3.185 15.555 3.185 15.555 3.46 15.325 3.46 15.325 3.185 13.85 3.185 13.85 3.83 12.565 3.83 12.565 3.185 10.555 3.185 10.555 3.83 10.325 3.83  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.385 4.59 2.385 3.58 2.615 3.58 2.615 4.59 6.865 4.59 6.865 3.58 7.095 3.58 7.095 4.59 13.87 4.59 20.875 4.59 20.875 4.15 21.105 4.15 21.105 4.59 25.355 4.59 25.355 3.875 25.585 3.875 25.585 4.59 27.775 4.59 27.875 4.59 28.56 4.59 28.56 5.49 27.875 5.49 27.775 5.49 13.87 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 28.56 -0.45 28.56 0.45 12.795 0.45 12.795 1.07 12.565 1.07 12.565 0.45 10.555 0.45 10.555 1.07 10.325 1.07 10.325 0.45 8.315 0.45 8.315 1.07 8.085 1.07 8.085 0.45 6.075 0.45 6.075 1.07 5.845 1.07 5.845 0.45 3.835 0.45 3.835 1.07 3.605 1.07 3.605 0.45 1.595 0.45 1.595 1.07 1.365 1.07 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.295 3.12 7.555 3.12 7.555 4.06 11.345 4.06 11.345 3.48 11.575 3.48 11.575 4.06 13.87 4.06 13.87 4.29 7.325 4.29 7.325 3.35 4.905 3.35 4.905 3.93 4.675 3.93 4.675 3.35 0.525 3.35 0.525 3.93 0.295 3.93  ;
        POLYGON 14.305 3.48 14.535 3.48 14.535 3.69 16.445 3.69 16.445 3.48 16.675 3.48 16.675 3.69 23.115 3.69 23.115 3.415 27.775 3.415 27.775 4.225 27.545 4.225 27.545 3.645 23.345 3.645 23.345 3.92 14.305 3.92  ;
        POLYGON 0.245 0.73 0.475 0.73 0.475 1.31 2.485 1.31 2.485 0.73 2.715 0.73 2.715 1.31 4.725 1.31 4.725 0.73 4.955 0.73 4.955 1.31 6.965 1.31 6.965 0.73 7.195 0.73 7.195 1.31 9.205 1.31 9.205 0.73 9.435 0.73 9.435 1.31 11.445 1.31 11.445 0.73 11.675 0.73 11.675 1.31 14.2 1.31 14.2 0.68 27.875 0.68 27.875 1.07 25.405 1.07 25.405 0.91 23.45 0.91 23.45 1.015 23.11 1.015 23.11 0.91 21.21 0.91 21.21 1.015 20.87 1.015 20.87 0.91 18.97 0.91 18.97 1.015 18.63 1.015 18.63 0.91 16.675 0.91 16.675 1.07 14.43 1.07 14.43 1.54 0.245 1.54  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai33_4
