# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.04 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.985 2.27 4.33 2.27 4.33 2.71 3.985 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.915 2.215 3.21 2.215 3.21 2.71 2.915 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.555 1.83 2.555  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.77 1.125 1.77 1.125 2.5 0.71 2.5  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.912 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.42 3.26 3.54 3.26 3.54 3.025 4.56 3.025 4.56 1.49 4.48 1.49 4.48 0.68 4.79 0.68 4.79 3.255 3.77 3.255 3.77 4.36 3.46 4.36 3.46 3.49 1.65 3.49 1.65 4.36 1.42 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.4 4.59 0.4 3.72 0.63 3.72 0.63 4.59 2.44 4.59 2.44 3.72 2.67 3.72 2.67 4.59 4.48 4.59 4.48 3.485 4.71 3.485 4.71 4.59 5.04 4.59 5.04 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 5.04 -0.45 5.04 0.45 0.63 0.45 0.63 1.49 0.4 1.49 0.4 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand4_1
