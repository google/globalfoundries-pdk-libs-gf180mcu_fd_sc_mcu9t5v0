# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 23.52 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 27.06 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.27 9.9 2.27 9.9 2.65 0.63 2.65  ;
        POLYGON 11.11 2.27 20.38 2.27 20.38 2.65 11.11 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 15.142 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 10.13 3.09 10.13 1.745 1.365 1.745 1.365 0.945 1.625 0.945 1.625 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 5.845 1.515 5.845 0.945 6.075 0.945 6.075 1.515 8.085 1.515 8.085 0.945 8.315 0.945 8.315 1.515 10.325 1.515 10.325 0.945 10.555 0.945 10.555 1.515 12.565 1.515 12.565 0.945 12.795 0.945 12.795 1.515 14.805 1.515 14.805 0.945 15.035 0.945 15.035 1.515 17.045 1.515 17.045 0.945 17.275 0.945 17.275 1.515 19.285 1.515 19.285 0.945 19.515 0.945 19.515 1.515 21.525 1.515 21.525 0.945 21.755 0.945 21.755 1.745 10.88 1.745 10.88 3.09 21.655 3.09 21.655 4.36 21.425 4.36 21.425 3.32 19.415 3.32 19.415 4.36 19.185 4.36 19.185 3.32 17.175 3.32 17.175 4.36 16.945 4.36 16.945 3.32 14.935 3.32 14.935 4.36 14.705 4.36 14.705 3.32 12.695 3.32 12.695 4.36 12.465 4.36 12.465 3.32 10.455 3.32 10.455 4.36 10.225 4.36 10.225 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.55 11.575 3.55 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 15.825 4.59 15.825 3.55 16.055 3.55 16.055 4.59 18.065 4.59 18.065 3.55 18.295 3.55 18.295 4.59 20.305 4.59 20.305 3.55 20.535 3.55 20.535 4.59 22.545 4.59 22.545 3.55 22.775 3.55 22.775 4.59 23.52 4.59 23.52 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 23.52 -0.45 23.52 0.45 22.875 0.45 22.875 1.285 22.645 1.285 22.645 0.45 20.635 0.45 20.635 1.285 20.405 1.285 20.405 0.45 18.395 0.45 18.395 1.285 18.165 1.285 18.165 0.45 16.155 0.45 16.155 1.285 15.925 1.285 15.925 0.45 13.915 0.45 13.915 1.285 13.685 1.285 13.685 0.45 11.675 0.45 11.675 1.285 11.445 1.285 11.445 0.45 9.435 0.45 9.435 1.285 9.205 1.285 9.205 0.45 7.195 0.45 7.195 1.285 6.965 1.285 6.965 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_20
