# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai31_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai31_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 7.59 2.27 7.99 2.27 7.99 1.77 10.39 1.77 10.39 2.27 11.1 2.27 11.1 2.5 10.16 2.5 10.16 2 8.25 2 8.25 2.5 7.59 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.355 2.215 5.585 2.215 5.585 2.73 9.59 2.73 9.59 2.27 9.93 2.27 9.93 2.73 13.005 2.73 13.005 2.215 13.235 2.215 13.235 2.96 5.355 2.96  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.27 1.77 1.53 1.77 1.53 2.27 3.89 2.27 3.89 2.5 1.27 2.5  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458 ;
    PORT
      LAYER METAL1 ;
        POLYGON 15.27 2.27 17.85 2.27 17.85 2.71 15.27 2.71  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.50965 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.96 3.605 11.395 3.605 11.395 3.19 13.465 3.19 13.465 1.985 10.62 1.985 10.62 1.54 7.825 1.54 7.825 1.605 1.695 1.605 1.695 1.54 1.365 1.54 1.365 1.14 1.86 1.14 1.86 1.375 3.55 1.375 3.55 1.14 3.89 1.14 3.89 1.375 5.19 1.375 5.19 1.14 6.13 1.14 6.13 1.375 7.66 1.375 7.66 1.14 8.37 1.14 8.37 1.31 10.27 1.31 10.27 1.14 10.85 1.14 10.85 1.755 12.565 1.755 12.565 1.14 12.795 1.14 12.795 1.755 13.695 1.755 13.695 3.09 17.745 3.09 17.745 4.36 17.515 4.36 17.515 3.32 15.555 3.32 15.555 4.36 15.325 4.36 15.325 3.42 11.625 3.42 11.625 3.89 6.96 3.89  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.55 1.595 3.55 1.595 4.59 3.555 4.59 3.555 3.55 3.785 3.55 3.785 4.59 13.87 4.59 14.305 4.59 14.305 3.875 14.535 3.875 14.535 4.59 16.495 4.59 16.495 3.55 16.725 3.55 16.725 4.59 18.635 4.59 18.635 3.55 18.865 3.55 18.865 4.59 18.915 4.59 19.6 4.59 19.6 5.49 18.915 5.49 13.87 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 19.6 -0.45 19.6 0.45 17.795 0.45 17.795 1.58 17.565 1.58 17.565 0.45 15.555 0.45 15.555 1.58 15.325 1.58 15.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 3.09 5.165 3.09 5.165 4.12 13.87 4.12 13.87 4.35 4.935 4.35 4.935 3.32 2.715 3.32 2.715 4.36 2.485 4.36 2.485 3.32 0.575 3.32 0.575 4.36 0.345 4.36  ;
        POLYGON 0.245 0.68 14.155 0.68 14.155 1.81 16.445 1.81 16.445 0.805 16.675 0.805 16.675 1.81 18.685 1.81 18.685 0.805 18.915 0.805 18.915 2.04 13.925 2.04 13.925 0.91 11.675 0.91 11.675 1.525 11.445 1.525 11.445 0.91 9.49 0.91 9.49 1.08 9.15 1.08 9.15 0.91 7.195 0.91 7.195 1.145 6.965 1.145 6.965 0.91 4.955 0.91 4.955 1.145 4.725 1.145 4.725 0.91 2.715 0.91 2.715 1.145 2.485 1.145 2.485 0.91 0.475 0.91 0.475 1.615 0.245 1.615  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai31_4
