# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__latq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.2 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.065 1.21 4.33 1.21 4.33 2.15 4.065 2.15  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.575 1.015 1.575 1.015 2.71 0.71 2.71  ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.605 0.68 9.93 0.68 9.93 4.08 9.605 4.08  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.27 1.595 3.27 1.595 4.59 2.315 4.59 3.485 4.59 3.485 3.27 3.715 3.27 3.715 4.59 7.465 4.59 7.465 3.27 7.695 3.27 7.695 4.59 9.115 4.59 10.625 4.59 10.625 3.27 10.855 3.27 10.855 4.59 11.2 4.59 11.2 5.49 9.115 5.49 2.315 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.2 -0.45 11.2 0.45 10.955 0.45 10.955 1.49 10.725 1.49 10.725 0.45 7.995 0.45 7.995 0.885 7.765 0.885 7.765 0.45 3.615 0.45 3.615 1.02 3.385 1.02 3.385 0.45 1.595 0.45 1.595 0.895 1.365 0.895 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 1.115 1.155 1.115 1.155 1.125 2.315 1.125 2.315 1.915 2.085 1.915 2.085 1.355 1.085 1.355 1.085 1.345 0.475 1.345 0.475 3.27 0.575 3.27 0.575 4.08 0.245 4.08  ;
        POLYGON 2.665 0.68 2.895 0.68 2.895 2.38 4.665 2.38 4.665 1.575 4.895 1.575 4.895 2.38 5.755 2.38 5.755 2.95 5.525 2.95 5.525 2.61 2.895 2.61 2.895 4.08 2.665 4.08  ;
        POLYGON 5.245 3.18 5.985 3.18 5.985 1.225 5.345 1.225 5.345 0.885 6.19 0.885 6.19 1.115 8.435 1.115 8.435 1.915 8.205 1.915 8.205 1.345 6.215 1.345 6.215 3.41 5.475 3.41 5.475 4.08 5.245 4.08  ;
        POLYGON 7.085 1.575 7.315 1.575 7.315 2.145 8.665 2.145 8.665 0.975 9.115 0.975 9.115 2.365 8.735 2.365 8.735 4.08 8.485 4.08 8.485 2.375 7.085 2.375  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latq_1
