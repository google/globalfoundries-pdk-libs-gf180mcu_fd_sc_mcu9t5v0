# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.4 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.88 2.33 2.09 2.33 2.09 2.715 0.88 2.715  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.125 2.285 5.465 2.285 5.465 2.71 5.125 2.71  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6224 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.705 0.84 7.13 0.84 7.13 3.72 6.705 3.72  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.375 4.59 1.375 3.845 1.605 3.845 1.605 4.59 5.685 4.59 5.685 3.88 5.915 3.88 5.915 4.59 6.355 4.59 6.41 4.59 7.725 4.59 7.725 3.88 7.955 3.88 7.955 4.59 8.4 4.59 8.4 5.49 6.41 5.49 6.355 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.4 -0.45 8.4 0.45 8.155 0.45 8.155 1.16 7.925 1.16 7.925 0.45 5.915 0.45 5.915 1.16 5.685 1.16 5.685 0.45 1.605 0.45 1.605 1.165 1.375 1.165 1.375 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.255 0.845 0.485 0.845 0.485 1.83 2.55 1.83 2.55 2.415 3.715 2.415 3.715 2.645 2.32 2.645 2.32 2.06 0.585 2.06 0.585 3.685 0.255 3.685  ;
        POLYGON 2.925 2.875 3.155 2.875 3.155 3.455 4.665 3.455 4.665 1.655 3.615 1.655 3.615 1.315 4.895 1.315 4.895 3.275 6.125 3.275 6.125 2.45 6.355 2.45 6.355 3.505 4.89 3.505 4.89 3.685 2.925 3.685  ;
        POLYGON 2.495 0.68 5.355 0.68 5.355 1.825 6.41 1.825 6.41 2.055 5.125 2.055 5.125 1.085 3.385 1.085 3.385 1.955 4.175 1.955 4.175 3.215 3.945 3.215 3.945 2.185 3.155 2.185 3.155 1.49 2.495 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_2
