# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 24.64 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.51 1.77 3.995 1.77 3.995 2.71 3.51 2.71  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 2.275 0.97 2.275 0.97 2.71 0.15 2.71  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER METAL1 ;
        POLYGON 18.63 1.77 19.425 1.77 19.425 2.71 18.63 2.71  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.27 2.275 2.09 2.275 2.09 2.71 1.27 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.31 2.275 7.13 2.275 7.13 2.71 6.31 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 23.67 0.845 24.285 0.845 24.285 4.06 23.67 4.06  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 3.4 1.545 3.4 1.545 4.59 5.145 4.59 5.145 3.25 5.375 3.25 5.375 4.59 7.45 4.59 7.45 3.97 7.79 3.97 7.79 4.59 9.675 4.59 10.17 4.59 12.595 4.59 12.595 3.835 12.825 3.835 12.825 4.59 14.955 4.59 14.955 3.09 15.185 3.09 15.185 4.59 16.865 4.59 18.955 4.59 18.955 3.4 19.185 3.4 19.185 4.59 20.205 4.59 21.195 4.59 21.195 4.31 21.425 4.31 21.425 4.59 22.985 4.59 22.985 3.25 23.215 3.25 23.215 4.59 23.44 4.59 24.64 4.59 24.64 5.49 23.44 5.49 20.205 5.49 16.865 5.49 10.17 5.49 9.675 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 24.64 -0.45 24.64 0.45 23.165 0.45 23.165 1.165 22.935 1.165 22.935 0.45 21.105 0.45 21.105 0.61 20.875 0.61 20.875 0.45 12.98 0.45 12.98 0.625 12.64 0.625 12.64 0.45 7.785 0.45 7.785 1.14 7.555 1.14 7.555 0.45 5.685 0.45 5.685 0.63 5.455 0.63 5.455 0.45 1.595 0.45 1.595 1.45 1.365 1.45 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.295 2.94 2.545 2.94 2.545 2.045 0.245 2.045 0.245 1.11 0.475 1.11 0.475 1.815 2.775 1.815 2.775 2.94 4.225 2.94 4.225 1.73 4.835 1.73 4.835 2.07 4.455 2.07 4.455 3.17 0.525 3.17 0.525 4.06 0.295 4.06  ;
        POLYGON 6.485 2.94 7.445 2.94 7.445 2.06 7.215 2.06 7.215 2.045 6.435 2.045 6.435 1.14 6.665 1.14 6.665 1.815 7.3 1.815 7.3 1.83 7.675 1.83 7.675 2.275 8.28 2.275 8.28 2.505 7.675 2.505 7.675 3.28 6.485 3.28  ;
        POLYGON 3.325 0.86 5.985 0.86 5.985 0.68 7.125 0.68 7.125 1.355 7.47 1.355 7.47 1.37 8.015 1.37 8.015 0.68 9.625 0.68 9.625 1.135 9.395 1.135 9.395 0.91 8.245 0.91 8.245 1.6 7.385 1.6 7.385 1.585 6.895 1.585 6.895 0.91 6.21 0.91 6.21 1.09 3.555 1.09 3.555 1.45 3.325 1.45  ;
        POLYGON 3.325 3.4 4.685 3.4 4.685 2.79 5.835 2.79 5.835 3.51 9.445 3.51 9.445 2.93 9.675 2.93 9.675 3.74 5.605 3.74 5.605 3.02 4.915 3.02 4.915 3.63 3.555 3.63 3.555 4.21 3.325 4.21  ;
        POLYGON 8.575 1.14 8.905 1.14 8.905 2.275 10.17 2.275 10.17 2.505 8.805 2.505 8.805 3.235 8.575 3.235  ;
        POLYGON 10.515 1.025 10.745 1.025 10.745 2.055 13.64 2.055 13.64 2.285 10.745 2.285 10.745 3.73 10.515 3.73  ;
        POLYGON 11.195 0.855 15.44 0.855 15.44 0.68 15.78 0.68 15.78 1.085 11.425 1.085 11.425 1.825 11.195 1.825  ;
        POLYGON 11.88 2.515 13.935 2.515 13.935 1.315 15.285 1.315 15.285 1.68 16.425 1.68 16.425 3.73 16.195 3.73 16.195 1.91 15.055 1.91 15.055 1.545 14.165 1.545 14.165 3.26 13.935 3.26 13.935 2.745 11.88 2.745  ;
        POLYGON 11.095 3.375 13.225 3.375 13.225 3.49 14.495 3.49 14.495 2.63 15.965 2.63 15.965 4.02 16.865 4.02 16.865 4.36 15.735 4.36 15.735 2.86 14.725 2.86 14.725 3.72 13.025 3.72 13.025 3.605 11.325 3.605 11.325 4.36 11.095 4.36  ;
        POLYGON 18.4 2.94 20.205 2.94 20.205 3.95 19.975 3.95 19.975 3.17 18.465 3.17 18.465 3.9 18.17 3.9 18.17 1.48 17.295 1.48 17.295 1.14 18.985 1.14 18.985 1.48 18.4 1.48  ;
        POLYGON 16.175 0.68 19.425 0.68 19.425 0.84 21.865 0.84 21.865 2.56 21.635 2.56 21.635 1.07 19.205 1.07 19.205 0.91 17.065 0.91 17.065 1.71 17.445 1.71 17.445 3.9 17.215 3.9 17.215 1.94 16.835 1.94 16.835 0.91 16.405 0.91 16.405 1.45 16.175 1.45  ;
        POLYGON 20.555 2.22 20.785 2.22 20.785 2.79 22.215 2.79 22.215 1.11 22.445 1.11 22.445 2.22 23.44 2.22 23.44 2.56 22.445 2.56 22.445 4.1 22.215 4.1 22.215 3.02 20.555 3.02  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1
