# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.242 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.13 2.27 5.64 2.27 5.64 2.65 0.13 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.926 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.135 2.84 12.91 2.84 13.5 2.84 13.5 2.04 8.135 2.04 8.135 0.68 8.365 0.68 8.365 1.755 10.375 1.755 10.375 0.68 10.605 0.68 10.605 1.755 12.385 1.755 12.385 0.68 12.845 0.68 12.845 1.755 14.855 1.755 14.855 0.68 15.085 0.68 15.085 1.755 17.095 1.755 17.095 0.68 17.325 0.68 17.325 1.755 19.335 1.755 19.335 0.68 19.565 0.68 19.565 1.985 14 1.985 14 2.84 19.465 2.84 19.465 4.36 19.235 4.36 19.235 3.32 17.225 3.32 17.225 4.36 16.995 4.36 16.995 3.32 14.985 3.32 14.985 4.36 14.755 4.36 14.755 3.32 12.91 3.32 12.745 3.32 12.745 4.36 12.515 4.36 12.515 3.32 10.505 3.32 10.505 4.36 10.275 4.36 10.275 3.32 8.365 3.32 8.365 4.36 8.135 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 2.435 4.59 2.435 3.55 2.665 3.55 2.665 4.59 4.675 4.59 4.675 3.55 4.905 3.55 4.905 4.59 6.915 4.59 6.915 3.55 7.145 3.55 7.145 4.59 9.155 4.59 9.155 3.875 9.385 3.875 9.385 4.59 11.395 4.59 11.395 3.55 11.625 3.55 11.625 4.59 12.91 4.59 13.635 4.59 13.635 3.55 13.865 3.55 13.865 4.59 15.875 4.59 15.875 3.55 16.105 3.55 16.105 4.59 18.115 4.59 18.115 3.55 18.345 3.55 18.345 4.59 19.63 4.59 20.355 4.59 20.355 3.55 20.585 3.55 20.585 4.59 21.28 4.59 21.28 5.49 19.63 5.49 12.91 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.685 0.45 20.685 1.49 20.455 1.49 20.455 0.45 18.445 0.45 18.445 1.49 18.215 1.49 18.215 0.45 16.205 0.45 16.205 1.49 15.975 1.49 15.975 0.45 13.965 0.45 13.965 1.49 13.735 1.49 13.735 0.45 11.725 0.45 11.725 1.49 11.495 1.49 11.495 0.45 9.485 0.45 9.485 1.49 9.255 1.49 9.255 0.45 7.245 0.45 7.245 1.49 7.015 1.49 7.015 0.45 5.005 0.45 5.005 1.49 4.775 1.49 4.775 0.45 2.765 0.45 2.765 1.49 2.535 1.49 2.535 0.45 0.525 0.45 0.525 1.49 0.295 1.49 0.295 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.415 2.88 5.895 2.88 5.895 2.04 1.415 2.04 1.415 0.68 1.645 0.68 1.645 1.72 3.655 1.72 3.655 0.68 3.885 0.68 3.885 1.72 5.895 1.72 5.895 0.68 6.225 0.68 6.225 2.27 12.91 2.27 12.91 2.5 6.225 2.5 6.225 4.36 5.82 4.36 5.82 3.32 3.785 3.32 3.785 4.36 3.555 4.36 3.555 3.32 1.645 3.32 1.645 4.36 1.415 4.36  ;
        POLYGON 14.23 2.215 19.63 2.215 19.63 2.555 14.23 2.555  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_12
