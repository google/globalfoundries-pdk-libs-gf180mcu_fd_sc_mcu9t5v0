# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.75 3.895 1.75 3.895 2.09 2.89 2.09  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.97 1.75 13.78 1.75 13.78 2.09 12.97 2.09  ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 2.33 1.57 2.33 1.57 2.71 0.15 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.37 2.875 19.365 2.875 19.595 2.875 19.595 1.625 17.37 1.625 17.37 0.815 17.6 0.815 17.6 1.395 19.61 1.395 19.61 0.815 19.84 0.815 19.84 3.685 19.41 3.685 19.41 3.215 19.365 3.215 17.605 3.215 17.605 3.685 17.37 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.105 4.59 3.105 3.09 3.335 3.09 3.335 4.59 4.795 4.59 7.185 4.59 7.185 3.56 7.415 3.56 7.415 4.59 8.435 4.59 8.925 4.59 8.925 3.39 9.155 3.39 9.155 4.59 9.65 4.59 10.225 4.59 13.33 4.59 13.33 4.345 13.56 4.345 13.56 4.59 15.06 4.59 15.37 4.59 15.37 3.875 15.605 3.875 15.605 4.59 16.345 4.59 16.345 3.875 16.58 3.875 16.58 4.59 18.39 4.59 18.39 3.875 18.62 3.875 18.62 4.585 19.365 4.585 20.43 4.585 20.43 3.875 20.66 3.875 20.66 4.59 21.28 4.59 21.28 5.49 19.365 5.49 15.06 5.49 10.225 5.49 9.65 5.49 8.435 5.49 4.795 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.96 0.45 20.96 1.165 20.73 1.165 20.73 0.45 18.72 0.45 18.72 1.165 18.49 1.165 18.49 0.45 16.535 0.45 16.535 0.64 13.34 0.64 13.34 1.37 13.11 1.37 13.11 0.45 8.535 0.45 8.535 1.37 8.305 1.37 8.305 0.45 3.455 0.45 3.455 1.37 3.225 1.37 3.225 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 1.685 0.245 1.685 0.245 1.315 0.475 1.315 0.475 1.455 2.035 1.455 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.125 1.26 4.575 1.26 4.575 3.73 4.125 3.73  ;
        POLYGON 2.615 2.63 3.895 2.63 3.895 4.02 4.795 4.02 4.795 4.36 3.665 4.36 3.665 2.86 2.615 2.86 2.615 3.685 2.385 3.685 2.385 1.26 2.715 1.26 2.715 1.6 2.615 1.6  ;
        POLYGON 6.165 3.09 8.435 3.09 8.435 3.9 8.205 3.9 8.205 3.32 6.395 3.32 6.395 3.9 6.165 3.9  ;
        POLYGON 5.375 2.63 9.65 2.63 9.65 2.86 5.375 2.86 5.375 3.73 5.145 3.73 5.145 1.26 5.695 1.26 5.695 1.6 5.375 1.6  ;
        POLYGON 6.69 2.06 9.75 2.06 9.75 1.26 9.98 1.26 9.98 2.2 10.225 2.2 10.225 4.03 9.995 4.03 9.995 2.43 9.765 2.43 9.765 2.29 6.69 2.29  ;
        POLYGON 6.145 1.6 9.29 1.6 9.29 0.8 11.685 0.8 11.685 3.1 11.455 3.1 11.455 1.03 10.64 1.03 10.64 2.06 10.41 2.06 10.41 1.03 9.52 1.03 9.52 1.83 6.375 1.83 6.375 2.06 6.145 2.06  ;
        POLYGON 11.99 1.26 12.265 1.26 12.265 3.56 11.99 3.56  ;
        POLYGON 10.87 1.26 11.1 1.26 11.1 3.22 11.245 3.22 11.245 3.8 14.83 3.8 14.83 2.415 15.06 2.415 15.06 4.03 10.87 4.03  ;
        POLYGON 12.67 2.76 14.35 2.76 14.35 1.955 15.53 1.955 15.53 1.315 15.76 1.315 15.76 1.955 19.365 1.955 19.365 2.185 14.58 2.185 14.58 3.215 12.67 3.215  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_4
