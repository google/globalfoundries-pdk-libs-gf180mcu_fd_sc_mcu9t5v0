# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi21_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.415 2.655 2.415 2.655 3.27 1.83 3.27  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.285 0.97 2.285 0.97 2.71 0.115 2.71  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.467 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.805 3.78 1.805 3.78 2.815 2.95 2.815  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 1.77 2.285 1.77 2.285 0.845 2.515 0.845 2.515 2.15 1.495 2.15 1.495 3.685 1.265 3.685  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.515 4.59 3.485 4.59 3.485 3.875 3.715 3.875 3.715 4.59 4.48 4.59 4.48 5.49 2.515 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 3.815 0.45 3.815 1.565 3.585 1.565 3.585 0.45 0.475 0.45 0.475 1.165 0.245 1.165 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.55 0.475 3.55 0.475 4.13 2.285 4.13 2.285 3.55 2.515 3.55 2.515 4.36 0.245 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi21_1
