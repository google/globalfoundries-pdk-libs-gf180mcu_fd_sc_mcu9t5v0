# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__or3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.72 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.27 1.07 2.27 1.07 2.71 0.71 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.795 2.215 2.09 2.215 2.09 2.71 1.795 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.545 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.915 2.215 3.21 2.215 3.21 2.71 2.915 2.71  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7295 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.63 2.89 4.905 2.89 4.905 0.68 5.135 0.68 5.135 4.36 4.63 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 3.555 4.59 3.555 3.55 3.785 3.55 3.785 4.59 4.505 4.59 5.925 4.59 5.925 3.55 6.155 3.55 6.155 4.59 6.72 4.59 6.72 5.49 4.505 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 6.72 -0.45 6.72 0.45 6.255 0.45 6.255 1.49 6.025 1.49 6.025 0.45 3.835 0.45 3.835 1.385 3.605 1.385 3.605 0.45 1.595 0.45 1.595 1.385 1.365 1.385 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 3.09 3.44 3.09 3.44 1.845 0.245 1.845 0.245 0.68 0.475 0.68 0.475 1.615 2.485 1.615 2.485 0.68 2.715 0.68 2.715 1.615 3.67 1.615 3.67 2.215 4.505 2.215 4.505 2.555 3.67 2.555 3.67 3.32 0.575 3.32 0.575 4.36 0.345 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or3_2
