* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__bufz_1 EN I Z VDD VNW VPW VSS
*.PININFO EN:I I:I Z:O VDD:P VNW:P VPW:P VSS:G
*.EQN Z=I
M_XX27 VSS EN NEN VPW nmos_5p0 W=0.590000U L=0.600000U
M_XX44 VSS NEN NI_N VPW nmos_5p0 W=0.590000U L=0.600000U
M_XX36 NI_N EN NI_P VPW nmos_5p0 W=0.590000U L=0.600000U
M_XX43 NI_N I VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_XX22 Z NI_N VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_XX28 VDD EN NEN VNW pmos_5p0 W=0.990000U L=0.500000U
M_XX45 NI_P EN VDD VNW pmos_5p0 W=0.990000U L=0.500000U
M_XX39 NI_N NEN NI_P VNW pmos_5p0 W=0.990000U L=0.500000U
M_XX46 NI_P I VDD VNW pmos_5p0 W=0.990000U L=0.500000U
M_XX21 VDD NI_P Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
