# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyc_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyc_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.2 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.77 0.97 1.77 0.97 2.56 0.63 2.56  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.23 2.89 10.295 2.89 10.69 2.89 10.69 0.68 10.92 0.68 10.92 4.36 10.59 4.36 10.59 3.27 10.295 3.27 10.23 3.27  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.84 4.59 4.44 4.59 8.44 4.59 10.295 4.59 11.2 4.59 11.2 5.49 10.295 5.49 8.44 5.49 4.44 5.49 0 5.49 0 4.59 1.61 4.59 1.61 3.88 4.44 3.88 8.44 3.88 9.02 3.88 9.02 4.22 8.44 4.22 4.44 4.22 1.84 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.2 -0.45 11.2 0.45 9.12 0.45 9.12 0.695 8.89 0.695 8.89 0.45 5.12 0.45 5.12 0.69 4.89 0.69 4.89 0.45 1.595 0.45 1.595 0.965 1.365 0.965 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.4 2.79 1.2 2.79 1.2 2.33 1.995 2.33 1.995 1.86 2.335 1.86 2.335 2.56 1.43 2.56 1.43 3.02 0.475 3.02 0.475 4.22 0.17 4.22 0.17 0.68 0.53 0.68 0.53 0.91 0.4 0.91  ;
        POLYGON 1.555 3.215 4.21 3.215 4.21 1.63 1.555 1.63 1.555 1.4 4.44 1.4 4.44 3.445 1.555 3.445  ;
        POLYGON 4.79 1.07 5.12 1.07 5.12 1.86 6.335 1.86 6.335 2.56 5.995 2.56 5.995 2.09 5.02 2.09 5.02 3.5 4.79 3.5  ;
        POLYGON 5.61 2.79 6.565 2.79 6.565 1.63 5.61 1.63 5.61 1.07 5.84 1.07 5.84 1.4 8.44 1.4 8.44 2.615 8.21 2.615 8.21 1.63 6.795 1.63 6.795 3.02 5.84 3.02 5.84 3.5 5.61 3.5  ;
        POLYGON 8.79 1.075 9.12 1.075 9.12 1.86 10.295 1.86 10.295 2.56 9.955 2.56 9.955 2.09 9.02 2.09 9.02 3.5 8.79 3.5  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyc_1
