# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8595 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.99 1.77 4.33 1.77 4.33 2.395 3.99 2.395 3.99 2 2.33 2 2.33 2.36 1.99 2.36  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8595 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.96 2.11 1.19 2.11 1.19 3.05 3.29 3.05 3.51 3.05 3.51 2.89 3.74 2.89 3.74 2.625 5.01 2.625 5.01 2.165 5.35 2.165 5.35 2.855 3.97 2.855 3.97 3.28 3.29 3.28 0.96 3.28  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.145 2.775 9.785 2.775 10.23 2.775 10.23 2.33 10.805 2.33 10.805 2.56 10.49 2.56 10.49 3.005 9.785 3.005 8.145 3.005  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.593 ;
    PORT
      LAYER METAL1 ;
        POLYGON 12.94 3.415 13.665 3.415 13.895 3.415 13.895 2 12.84 2 12.84 0.845 13.07 0.845 13.07 1.77 15.08 1.77 15.08 0.845 15.31 0.845 15.31 1.885 17.32 1.885 17.32 0.845 17.55 0.845 17.55 4.345 17.22 4.345 17.22 2.115 15.26 2.115 15.26 4.345 15.03 4.345 15.03 2.15 14.125 2.15 14.125 3.645 13.665 3.645 13.17 3.645 13.17 4.345 12.94 4.345  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 2.385 4.59 2.385 3.535 2.615 3.535 2.615 4.59 3.29 4.59 6.11 4.59 8.64 4.59 8.64 3.535 8.87 3.535 8.87 4.59 9.785 4.59 12.35 4.59 13.665 4.59 13.96 4.59 13.96 3.875 14.19 3.875 14.19 4.59 16.15 4.59 16.15 3.875 16.38 3.875 16.38 4.59 17.92 4.59 17.92 5.49 13.665 5.49 12.35 5.49 9.785 5.49 6.11 5.49 3.29 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 16.43 0.45 16.43 1.655 16.2 1.655 16.2 0.45 14.19 0.45 14.19 1.165 13.96 1.165 13.96 0.45 12.35 0.45 12.35 1.165 12.12 1.165 12.12 0.45 9.19 0.45 9.19 1.165 8.96 1.165 8.96 0.45 5.645 0.45 5.645 0.845 6.73 0.845 6.73 1.48 6.5 1.48 6.5 1.185 5.415 1.185 5.415 0.45 2.715 0.45 2.715 1.185 2.485 1.185 2.485 0.45 0.475 0.45 0.475 1.185 0.245 1.185 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 1.65 1.365 1.65 1.365 0.845 1.65 0.845 1.65 2.59 3.29 2.59 3.29 2.82 1.42 2.82 1.42 1.88 0.575 1.88 0.575 3.875 0.345 3.875  ;
        POLYGON 3.605 3.535 3.835 3.535 3.835 4.105 5.88 4.105 5.88 3.535 6.11 3.535 6.11 4.335 3.605 4.335  ;
        POLYGON 6.6 2.68 7.62 2.68 7.62 1.14 7.85 1.14 7.85 2.315 9.785 2.315 9.785 2.545 7.85 2.545 7.85 2.91 6.83 2.91 6.83 3.875 6.6 3.875  ;
        POLYGON 4.625 3.085 5.58 3.085 5.58 1.935 4.56 1.935 4.56 1.13 3.55 1.13 3.55 0.9 4.79 0.9 4.79 1.705 5.63 1.705 5.63 1.71 7.04 1.71 7.04 0.68 8.31 0.68 8.31 1.855 11.825 1.855 11.825 2.085 8.08 2.085 8.08 0.91 7.27 0.91 7.27 2.45 7.04 2.45 7.04 1.94 5.81 1.94 5.81 3.315 4.855 3.315 4.855 3.875 4.625 3.875  ;
        POLYGON 10.08 3.55 10.31 3.55 10.31 4.13 12.12 4.13 12.12 3.55 12.35 3.55 12.35 4.36 10.08 4.36  ;
        POLYGON 11.1 2.315 12.055 2.315 12.055 1.625 10.08 1.625 10.08 0.815 10.31 0.815 10.31 1.395 12.285 1.395 12.285 2.23 13.665 2.23 13.665 2.545 11.33 2.545 11.33 3.9 11.1 3.9  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_4
