* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__or4_4 A1 A2 A3 A4 Z VDD VNW VPW VSS
*.PININFO A1:I A2:I A3:I A4:I Z:O VDD:P VNW:P VPW:P VSS:G
*.EQN Z=(((A1 + A2) + A3) + A4)
M_i_5_1_x2_1 Z_neg A4 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_4_1_x2_1 VSS A3 Z_neg VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3_1_x2_1 Z_neg A2 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_1_x2_1 VSS A1 Z_neg VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_2_1_x2_0 Z_neg A1 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_3_1_x2_0 VSS A2 Z_neg VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_4_1_x2_0 Z_neg A3 VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_5_1_x2_0 VSS A4 Z_neg VPW nmos_5p0 W=0.790000U L=0.600000U
M_i_0_3_x4_3 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3_x4_2 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3_x4_1 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3_x4_0 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9_0_m2_1 net_2_0_1 A4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0_m2_1 net_1_0_1 A3 net_2_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0_m2_1 net_0_0_1 A2 net_1_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0_m2_1 Z_neg A1 net_0_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6_0_m2_0 net_0_0_0 A1 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0_m2_0 net_1_0_0 A2 net_0_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_8_0_m2_0 net_2_0_0 A3 net_1_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_9_0_m2_0 VDD A4 net_2_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3_x4_3 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3_x4_2 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3_x4_1 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_3_x4_0 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
