# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.28 2.33 3.915 2.33 3.915 2.71 3.28 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.83 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.865 1.66 14.15 1.66 14.15 1.21 15.07 1.21 15.07 1.59 14.38 1.59 14.38 2 13.865 2  ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 2.15 0.97 2.15 0.97 2.71 0.66 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.325 0.845 16.65 0.845 16.65 3.685 16.345 3.685 16.345 2.19 16.325 2.19  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.285 4.59 1.285 3.425 1.515 3.425 1.515 4.59 2.01 4.59 3.245 4.59 3.245 3.615 3.475 3.615 3.475 4.59 4.99 4.59 7.325 4.59 7.325 3.615 7.555 3.615 7.555 4.59 8.575 4.59 9.065 4.59 9.065 3.33 9.295 3.33 9.295 4.59 9.79 4.59 10.315 4.59 13.365 4.59 13.365 4.19 13.595 4.19 13.595 4.59 15.295 4.59 15.625 4.59 15.625 3.31 15.855 3.31 15.855 4.59 16.1 4.59 17.365 4.59 17.365 3.875 17.595 3.875 17.595 4.59 17.92 4.59 17.92 5.49 16.1 5.49 15.295 5.49 10.315 5.49 9.79 5.49 8.575 5.49 4.99 5.49 2.01 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 17.675 0.45 17.675 1.165 17.445 1.165 17.445 0.45 13.415 0.45 13.415 1.2 13.185 1.2 13.185 0.45 8.935 0.45 8.935 1.2 8.705 1.2 8.705 0.45 3.455 0.45 3.455 1.2 3.225 1.2 3.225 0.45 1.615 0.45 1.615 1.225 1.385 1.225 1.385 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.265 2.875 0.495 2.875 0.495 2.94 1.2 2.94 1.2 1.685 0.21 1.685 0.21 1.37 1.085 1.37 1.085 1.455 1.43 1.455 1.43 2.03 2.01 2.03 2.01 2.26 1.43 2.26 1.43 3.17 0.495 3.17 0.495 3.685 0.265 3.685  ;
        POLYGON 4.265 1.2 4.575 1.2 4.575 3.785 4.265 3.785  ;
        POLYGON 2.305 1.315 2.735 1.315 2.735 3.155 3.935 3.155 3.935 4.13 4.99 4.13 4.99 4.36 3.705 4.36 3.705 3.385 2.535 3.385 2.535 3.685 2.305 3.685  ;
        POLYGON 6.305 3.145 8.575 3.145 8.575 3.955 8.345 3.955 8.345 3.375 6.535 3.375 6.535 3.955 6.305 3.955  ;
        POLYGON 5.52 2.685 9.79 2.685 9.79 2.915 5.515 2.915 5.515 3.785 5.285 3.785 5.285 1.2 5.695 1.2 5.695 1.54 5.52 1.54  ;
        POLYGON 6.83 2.175 9.825 2.175 9.825 1.2 10.055 1.2 10.055 2.23 10.315 2.23 10.315 3.97 10.085 3.97 10.085 2.46 9.855 2.46 9.855 2.405 6.83 2.405  ;
        POLYGON 5.85 1.715 9.365 1.715 9.365 0.74 11.83 0.74 11.83 2.985 11.485 2.985 11.485 0.97 10.515 0.97 10.515 2 10.285 2 10.285 0.97 9.595 0.97 9.595 1.945 5.85 1.945  ;
        POLYGON 12.065 1.2 12.355 1.2 12.355 3.5 12.065 3.5  ;
        POLYGON 10.945 1.2 11.175 1.2 11.175 3.16 11.335 3.16 11.335 3.73 15.065 3.73 15.065 2.7 15.295 2.7 15.295 3.96 11.335 3.96 11.335 3.97 10.945 3.97  ;
        POLYGON 12.65 2.24 15.605 2.24 15.605 1.29 15.835 1.29 15.835 2.24 16.1 2.24 16.1 2.47 14.835 2.47 14.835 3.5 14.605 3.5 14.605 2.65 12.65 2.65  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_1
