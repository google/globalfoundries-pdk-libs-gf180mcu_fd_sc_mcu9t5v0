# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi221_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 22.4 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.21 1.91 16.95 1.91 16.95 1.21 18.23 1.21 18.23 1.72 19.77 1.72 19.77 2.37 21.45 2.37 21.45 2.6 19.54 2.6 19.54 1.95 18 1.95 18 1.44 17.27 1.44 17.27 2.4 16.93 2.4 16.93 2.14 14.55 2.14 14.55 2.5 14.21 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.15 2.37 16.7 2.37 16.7 2.63 17.51 2.63 17.51 1.77 17.77 1.77 17.77 2.27 19.31 2.27 19.31 2.5 17.74 2.5 17.74 2.86 16.47 2.86 16.47 2.6 16.15 2.6  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.7 1.855 3.51 1.855 3.51 1.21 3.77 1.21 3.77 1.755 6.425 1.755 6.425 2.37 8.16 2.37 8.16 2.6 6.195 2.6 6.195 1.985 3.925 1.985 3.925 2.4 3.695 2.4 3.695 2.085 1.04 2.085 1.04 2.6 0.7 2.6  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.504 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 2.315 1.985 2.315 1.985 2.63 5.735 2.63 5.735 2.215 5.965 2.215 5.965 2.86 1.27 2.86  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.11 2.27 9.65 2.27 9.65 2.71 9.11 2.71  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.0645 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 1.395 3.05 1.395 3.05 0.735 4.66 0.735 4.66 1.25 8.555 1.25 8.555 0.68 8.785 0.68 8.785 1.25 11.165 1.25 11.165 0.68 11.395 0.68 11.395 1.25 13.405 1.25 13.405 0.68 13.635 0.68 13.635 1.25 16.49 1.25 16.49 0.735 18.69 0.735 18.69 1.26 21.745 1.26 21.745 0.68 21.975 0.68 21.975 1.49 18.46 1.49 18.46 0.965 16.72 0.965 16.72 1.48 13.85 1.48 13.85 3.09 20.955 3.09 20.955 3.9 20.725 3.9 20.725 3.32 18.915 3.32 18.915 3.9 18.685 3.9 18.685 3.32 16.875 3.32 16.875 3.9 16.645 3.9 16.645 3.32 14.835 3.32 14.835 3.9 14.605 3.9 14.605 3.32 13.59 3.32 13.59 1.48 4.43 1.48 4.43 0.965 3.28 0.965 3.28 1.625 0.245 1.625  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.09 0.525 3.09 0.525 4.59 2.335 4.59 2.335 3.55 2.565 3.55 2.565 4.59 4.375 4.59 4.375 3.55 4.605 3.55 4.605 4.59 6.415 4.59 6.415 3.55 6.645 3.55 6.645 4.59 8.455 4.59 8.455 3.55 8.685 3.55 8.685 4.59 21.975 4.59 22.4 4.59 22.4 5.49 21.975 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 22.4 -0.45 22.4 0.45 19.935 0.45 19.935 1.02 19.705 1.02 19.705 0.45 15.855 0.45 15.855 1.02 15.625 1.02 15.625 0.45 12.515 0.45 12.515 1.02 12.285 1.02 12.285 0.45 10.275 0.45 10.275 1.02 10.045 1.02 10.045 0.45 6.645 0.45 6.645 1.02 6.415 1.02 6.415 0.45 2.565 0.45 2.565 1.165 2.335 1.165 2.335 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.315 3.09 10.34 3.09 10.34 3.075 12.465 3.075 12.465 3.9 12.235 3.9 12.235 3.305 10.425 3.305 10.425 3.9 10.195 3.9 10.195 3.32 7.665 3.32 7.665 3.9 7.435 3.9 7.435 3.32 5.625 3.32 5.625 3.9 5.395 3.9 5.395 3.32 3.585 3.32 3.585 3.9 3.355 3.9 3.355 3.32 1.545 3.32 1.545 3.9 1.315 3.9  ;
        POLYGON 9.175 3.55 9.405 3.55 9.405 4.13 11.215 4.13 11.215 3.535 11.445 3.535 11.445 4.13 13.305 4.13 13.305 3.545 13.535 3.545 13.535 4.13 15.625 4.13 15.625 3.55 15.855 3.55 15.855 4.13 17.665 4.13 17.665 3.55 17.895 3.55 17.895 4.13 19.705 4.13 19.705 3.55 19.935 3.55 19.935 4.13 21.745 4.13 21.745 3.09 21.975 3.09 21.975 4.36 9.175 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi221_4
