# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.72 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.075 1.77 3.975 1.77 3.975 2.15 3.075 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.435 1.21 14.97 1.21 14.97 1.59 14.665 1.59 14.665 2.115 14.435 2.115  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.24 1.39 2.24 1.39 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER METAL1 ;
        POLYGON 19.125 0.845 19.45 0.845 19.45 3.685 19.125 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.895 1.595 3.895 1.595 4.59 2.035 4.59 3.305 4.59 3.305 3.615 3.535 3.615 3.535 4.59 5.295 4.59 7.475 4.59 7.475 3.615 7.705 3.615 7.705 4.59 9.875 4.59 9.875 3.83 10.105 3.83 10.105 4.59 11.445 4.59 13.855 4.59 13.855 3.515 14.085 3.515 14.085 4.59 15.105 4.59 15.895 4.59 15.895 3.045 16.125 3.045 16.125 4.59 18.105 4.59 18.105 3.875 18.335 3.875 18.335 4.59 18.775 4.59 20.145 4.59 20.145 3.875 20.375 3.875 20.375 4.59 20.72 4.59 20.72 5.49 18.775 5.49 15.105 5.49 11.445 5.49 5.295 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 20.72 -0.45 20.72 0.45 20.475 0.45 20.475 1.165 20.245 1.165 20.245 0.45 18.235 0.45 18.235 1.165 18.005 1.165 18.005 0.45 16.345 0.45 16.345 1.165 16.115 1.165 16.115 0.45 7.705 0.45 7.705 1.32 7.475 1.32 7.475 0.45 3.435 0.45 3.435 1.32 3.205 1.32 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 2.9 0.575 2.9 0.575 3.01 1.805 3.01 1.805 1.74 0.245 1.74 0.245 1.315 0.475 1.315 0.475 1.51 2.035 1.51 2.035 3.24 0.345 3.24  ;
        POLYGON 4.325 1.21 4.555 1.21 4.555 3.785 4.325 3.785  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 2.985 3.995 2.985 3.995 4.13 5.295 4.13 5.295 4.36 3.765 4.36 3.765 3.215 2.385 3.215  ;
        POLYGON 5.445 1.21 5.675 1.21 5.675 2.185 6.64 2.185 6.64 2.11 8.42 2.11 8.42 2.34 6.81 2.34 6.81 2.415 5.82 2.415 5.82 3.785 5.445 3.785  ;
        POLYGON 6.13 1.65 7.935 1.65 7.935 0.68 10.38 0.68 10.38 0.91 8.165 0.91 8.165 1.88 6.47 1.88 6.47 1.955 6.13 1.955  ;
        POLYGON 6.98 2.57 9.655 2.57 9.655 1.315 9.885 1.315 9.885 2.57 11.005 2.57 11.005 3.215 10.775 3.215 10.775 2.8 8.805 2.8 8.805 3.315 8.575 3.315 8.575 2.8 6.98 2.8  ;
        POLYGON 6.115 3.155 8.165 3.155 8.165 3.545 9.425 3.545 9.425 3.37 10.445 3.37 10.445 3.445 11.445 3.445 11.445 4.315 11.215 4.315 11.215 3.675 10.275 3.675 10.275 3.6 9.65 3.6 9.65 3.775 7.935 3.775 7.935 3.385 6.455 3.385 6.455 4.36 6.115 4.36  ;
        POLYGON 13.365 2.985 15.105 2.985 15.105 3.795 14.875 3.795 14.875 3.215 13.135 3.215 13.135 1.655 11.895 1.655 11.895 1.21 14.165 1.21 14.165 1.55 13.365 1.55  ;
        POLYGON 10.775 0.75 15.43 0.75 15.43 1.83 16.84 1.83 16.84 2.06 15.2 2.06 15.2 0.98 11.665 0.98 11.665 1.885 12.025 1.885 12.025 3.685 11.795 3.685 11.795 2.115 11.435 2.115 11.435 0.98 11.005 0.98 11.005 1.425 10.775 1.425  ;
        POLYGON 15.455 2.29 17.215 2.29 17.215 0.845 17.465 0.845 17.465 1.775 18.775 1.775 18.775 2.115 17.445 2.115 17.445 3.685 17.135 3.685 17.135 2.63 15.455 2.63  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_2
