# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi22_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.36 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.21 2.27 11.66 2.27 11.66 2.63 14.185 2.63 14.185 2.215 14.415 2.215 14.415 2.86 11.44 2.86 11.44 2.71 11.21 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.325 1.77 13.185 1.77 13.185 0.68 16.355 0.68 16.355 2.555 16.125 2.555 16.125 0.91 13.415 0.91 13.415 2.4 12.47 2.4 12.47 2 9.555 2 9.555 2.555 9.325 2.555  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.81 2.27 3.21 2.27 3.21 2.785 4.205 2.785 4.205 2.27 6.07 2.27 6.07 2.5 4.435 2.5 4.435 3.015 2.81 3.015  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 1.77 7.715 1.77 7.715 2.215 7.955 2.215 7.955 2.555 7.485 2.555 7.485 2 3.975 2 3.975 2.555 3.745 2.555 3.745 2 0.915 2 0.915 2.555 0.15 2.555  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.552 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.095 3.08 11.245 3.08 11.245 3.09 14.765 3.09 14.765 1.14 14.995 1.14 14.995 3.09 16.015 3.09 16.015 3.9 15.27 3.9 15.27 3.32 13.975 3.32 13.975 3.9 13.745 3.9 13.745 3.32 11.935 3.32 11.935 3.9 11.705 3.9 11.705 3.32 11.195 3.32 11.195 3.315 10.965 3.315 10.965 3.31 9.895 3.31 9.895 3.9 8.865 3.9 8.865 1.985 7.945 1.985 7.945 1.54 2.285 1.54 2.285 0.73 2.515 0.73 2.515 1.31 6.365 1.31 6.365 0.73 6.595 0.73 6.595 1.31 8.175 1.31 8.175 1.755 8.865 1.755 8.865 0.73 10.915 0.73 10.915 1.54 9.095 1.54  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.245 1.495 3.245 1.495 4.59 3.305 4.59 3.305 3.705 3.535 3.705 3.535 4.59 5.345 4.59 5.345 3.705 5.575 3.705 5.575 4.59 7.385 4.59 7.385 3.705 7.615 3.705 7.615 4.59 17.035 4.59 17.36 4.59 17.36 5.49 17.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 17.36 -0.45 17.36 0.45 17.035 0.45 17.035 1.54 16.805 1.54 16.805 0.45 12.955 0.45 12.955 1.54 12.725 1.54 12.725 0.45 8.635 0.45 8.635 1.525 8.405 1.525 8.405 0.45 4.555 0.45 4.555 1.07 4.325 1.07 4.325 0.45 0.475 0.45 0.475 1.54 0.245 1.54 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 2.785 2.38 2.785 2.38 3.245 8.635 3.245 8.635 4.13 10.685 4.13 10.685 3.54 10.915 3.54 10.915 4.13 12.725 4.13 12.725 3.55 12.955 3.55 12.955 4.13 14.765 4.13 14.765 3.55 14.995 3.55 14.995 4.13 16.805 4.13 16.805 3.245 17.035 3.245 17.035 4.36 8.405 4.36 8.405 3.475 6.595 3.475 6.595 4.055 6.365 4.055 6.365 3.475 4.555 3.475 4.555 4.055 4.325 4.055 4.325 3.475 2.515 3.475 2.515 4.055 2.15 4.055 2.15 3.015 0.475 3.015 0.475 4.055 0.245 4.055  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi22_4
