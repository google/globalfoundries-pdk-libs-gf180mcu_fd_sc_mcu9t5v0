# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.02 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 2.275 3.81 2.275 3.81 2.505 3.21 2.505 3.21 3.27 2.95 3.27  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.322 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.925 1.76 6.115 1.76 6.115 2.56 5.885 2.56 5.885 1.99 4.755 1.99 4.755 2.71 4.07 2.71 4.07 1.99 1.155 1.99 1.155 2.56 0.925 2.56  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.44 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.275 2.65 2.275 2.65 2.71 1.83 2.71  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.302 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.11 1.77 9.535 1.77 9.535 2.71 9.11 2.71  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.47 1.21 12.945 1.21 12.945 0.79 13.175 0.79 13.175 4.31 12.945 4.31 12.945 2.15 12.47 2.15  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.88 1.595 3.88 1.595 4.59 3.425 4.59 3.425 4.42 3.655 4.42 3.655 4.59 7.565 4.59 7.565 3.5 7.795 3.5 7.795 4.59 8.235 4.59 9.985 4.59 9.985 3.88 10.215 3.88 10.215 4.59 11.825 4.59 11.825 3.88 12.055 3.88 12.055 4.59 12.24 4.59 14.065 4.59 14.065 3.88 14.295 3.88 14.295 4.59 14.56 4.59 14.56 5.49 12.24 5.49 8.235 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 14.295 0.45 14.295 1.6 14.065 1.6 14.065 0.45 12.055 0.45 12.055 1.53 11.825 1.53 11.825 0.45 7.835 0.45 7.835 1.13 7.605 1.13 7.605 0.45 1.815 0.45 1.815 1.13 1.585 1.13 1.585 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.79 0.695 0.79 0.695 3.42 2.665 3.42 2.665 3.5 5.125 3.5 5.125 2.22 5.355 2.22 5.355 3.73 2.49 3.73 2.49 3.65 0.475 3.65 0.475 4.31 0.245 4.31  ;
        POLYGON 2.085 3.88 2.315 3.88 2.315 3.96 5.605 3.96 5.605 2.79 6.345 2.79 6.345 1.13 4.805 1.13 4.805 0.79 6.575 0.79 6.575 2.79 8.005 2.79 8.005 2.22 8.235 2.22 8.235 3.02 5.835 3.02 5.835 4.31 5.605 4.31 5.605 4.19 2.315 4.19 2.315 4.22 2.085 4.22  ;
        POLYGON 8.865 3.42 9.765 3.42 9.765 1.54 8.21 1.54 8.21 1.99 7.365 1.99 7.365 2.56 7.135 2.56 7.135 1.76 7.98 1.76 7.98 1.31 9.745 1.31 9.745 0.79 9.995 0.79 9.995 2.22 11.375 2.22 11.375 2.56 9.995 2.56 9.995 3.65 9.095 3.65 9.095 4.31 8.865 4.31  ;
        POLYGON 10.705 3.42 12.01 3.42 12.01 1.99 10.705 1.99 10.705 0.79 10.935 0.79 10.935 1.76 12.24 1.76 12.24 3.65 10.935 3.65 10.935 4.31 10.705 4.31  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_2
