* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2 D RN SE SI CLK Q VDD VNW VPW VSS
*.PININFO D:I RN:I SE:I SI:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G
M_tn17 net3 SE VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn7 VSS SI net13 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn6 net13 SE net10 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn11 net10 D net5 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn16 net5 net3 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn10 ncki CLK VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn13 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn15 net10 ncki net1 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn14 net1 cki net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn8 net12 net2 net15 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn9 VSS RN net12 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn18 VSS net1 net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn0 net8 cki net2 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn1 net11 ncki net8 VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn12 net11 net4 VSS VPW nmos_5p0 W=0.590000U L=0.600000U
M_tn5 net0 RN VSS VPW nmos_5p0 W=1.000000U L=0.600000U
M_tn4 net4 net8 net0 VPW nmos_5p0 W=1.000000U L=0.600000U
M_tn3_17 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp17 net3 SE VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp16 net7 SI VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp13 net6 net3 net7 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp9 net14 D net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp14 VDD SE net14 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp8 ncki CLK VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp11 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp15 net1 cki net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net9 ncki net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 VDD net2 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net9 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 VDD net1 net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net2 ncki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 cki net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 RN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp4 VDD net8 net4 VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp1_16 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
