# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.475 2.215 3.77 2.215 3.77 2.71 3.475 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.215 2.135 2.215 2.135 2.94 5.215 2.94 5.215 2.215 5.445 2.215 5.445 3.17 1.83 3.17  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.215 1.495 2.215 1.495 3.4 6.31 3.4 6.31 2.215 6.57 2.215 6.57 3.63 1.265 3.63  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.6514 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 1.21 2.485 1.21 2.485 0.68 2.715 0.68 2.715 1.25 4.725 1.25 4.725 0.68 4.955 0.68 4.955 1.25 6.965 1.25 6.965 0.68 7.195 0.68 7.195 1.48 1.035 1.48 1.035 3.93 3.84 3.93 3.84 4.16 0.805 4.16 0.805 1.59 0.245 1.59  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.875 0.575 3.875 0.575 4.59 6.865 4.59 6.865 3.875 7.095 3.875 7.095 4.59 7.84 4.59 7.84 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 6.075 0.45 6.075 1.02 5.845 1.02 5.845 0.45 3.835 0.45 3.835 1.02 3.605 1.02 3.605 0.45 1.595 0.45 1.595 0.98 1.365 0.98 1.365 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor3_2
