# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nand2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.04 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.685 1.83 2.715 1.83 2.715 2.305 1.685 2.305  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.21 0.97 1.21 0.97 2.94 3.015 2.94 3.015 1.83 4.03 1.83 4.03 2.1 3.245 2.1 3.245 3.17 0.71 3.17  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3972 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.265 3.4 3.39 3.4 3.39 3.35 4.07 3.35 4.07 2.33 4.26 2.33 4.26 1.59 2.285 1.59 2.285 0.68 2.515 0.68 2.515 1.21 4.49 1.21 4.49 3.58 3.535 3.58 3.535 4.21 3.305 4.21 3.305 3.63 1.495 3.63 1.495 4.21 1.265 4.21  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.86 0.475 3.86 0.475 4.59 2.285 4.59 2.285 3.86 2.515 3.86 2.515 4.59 4.325 4.59 4.325 3.86 4.555 3.86 4.555 4.59 5.04 4.59 5.04 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 5.04 -0.45 5.04 0.45 4.555 0.45 4.555 0.695 4.325 0.695 4.325 0.45 0.475 0.45 0.475 1.165 0.245 1.165 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand2_2
