# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi222_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.7 2.345 11.775 2.345 11.775 1.21 12.96 1.21 12.96 2.575 9.7 2.575  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.945 1.21 11.05 1.21 11.05 2.115 9.945 2.115  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.605 2.38 7.605 2.38 7.605 1.77 8.81 1.77 8.81 2.61 5.605 2.61  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.255 1.77 6.77 1.77 6.77 2.15 5.255 2.15  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 2.415 4.065 2.415 4.065 2.645 0.97 2.645 0.97 3.27 0.115 3.27  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.77 2.09 1.77 2.09 2.15 0.825 2.15  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.2758 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 0.68 0.51 0.68 0.51 0.925 4.98 0.925 4.98 0.68 5.21 0.68 5.21 0.925 9.16 0.925 9.16 0.845 9.47 0.845 9.47 2.875 13.255 2.875 13.255 0.845 13.485 0.845 13.485 3.105 12.465 3.105 12.465 3.685 12.235 3.685 12.235 3.105 10.425 3.105 10.425 3.685 10.195 3.685 10.195 3.105 9.04 3.105 9.04 1.49 0.28 1.49 0.28 1.01 0.28 0.925  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.28 4.59 0.28 3.875 0.51 3.875 0.51 4.59 2.32 4.59 2.32 3.875 2.55 3.875 2.55 4.59 4.36 4.59 4.36 3.875 4.59 3.875 4.59 4.59 13.485 4.59 14 4.59 14 5.49 13.485 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14 -0.45 14 0.45 11.445 0.45 11.445 0.695 11.215 0.695 11.215 0.45 7.35 0.45 7.35 0.695 7.12 0.695 7.12 0.45 2.55 0.45 2.55 0.695 2.32 0.695 2.32 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.3 2.875 8.37 2.875 8.37 3.685 8.14 3.685 8.14 3.105 6.33 3.105 6.33 3.685 6.1 3.685 6.1 3.105 3.57 3.105 3.57 3.685 3.34 3.685 3.34 3.105 1.53 3.105 1.53 3.685 1.3 3.685  ;
        POLYGON 5.08 3.335 5.31 3.335 5.31 3.915 7.12 3.915 7.12 3.335 7.35 3.335 7.35 3.915 9.16 3.915 9.16 3.335 9.39 3.335 9.39 3.915 11.215 3.915 11.215 3.335 11.445 3.335 11.445 3.915 13.255 3.915 13.255 3.335 13.485 3.335 13.485 4.145 5.08 4.145  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi222_2
