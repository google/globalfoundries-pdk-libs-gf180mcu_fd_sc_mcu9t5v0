# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.945 2.31 3.77 2.31 3.77 2.71 2.945 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.03 ;
    PORT
      LAYER METAL1 ;
        POLYGON 13.59 1.21 13.91 1.21 13.91 2.025 13.59 2.025  ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.665 2.235 1.575 2.235 1.575 2.71 0.665 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 15.83 3.45 15.93 3.45 16.16 3.45 16.16 0.845 16.39 0.845 16.39 3.83 15.93 3.83 15.83 3.83  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.305 4.59 1.305 3.425 1.535 3.425 1.535 4.59 2.035 4.59 3.045 4.59 3.045 3.515 3.275 3.515 3.275 4.59 5.755 4.59 7.125 4.59 7.125 3.515 7.355 3.515 7.355 4.59 8.375 4.59 8.865 4.59 8.865 3.355 9.095 3.355 9.095 4.59 9.59 4.59 10.115 4.59 13.185 4.59 13.185 4.26 13.525 4.26 13.525 4.59 14.95 4.59 15.28 4.59 15.28 3.735 15.51 3.735 15.51 4.59 15.93 4.59 17.18 4.59 17.18 3.875 17.41 3.875 17.41 4.59 17.92 4.59 17.92 5.49 15.93 5.49 14.95 5.49 10.115 5.49 9.59 5.49 8.375 5.49 5.755 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 17.51 0.45 17.51 1.165 17.28 1.165 17.28 0.45 13.25 0.45 13.25 1.225 13.02 1.225 13.02 0.45 8.475 0.45 8.475 1.225 8.245 1.225 8.245 0.45 3.435 0.45 3.435 1.225 3.205 1.225 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.285 2.94 1.805 2.94 1.805 1.74 0.245 1.74 0.245 1.315 0.475 1.315 0.475 1.51 2.035 1.51 2.035 3.17 0.515 3.17 0.515 3.75 0.285 3.75  ;
        POLYGON 4.065 1.28 4.61 1.28 4.61 1.51 4.295 1.51 4.295 3.685 4.065 3.685  ;
        POLYGON 2.325 1.315 2.715 1.315 2.715 3.055 3.735 3.055 3.735 3.975 5.755 3.975 5.755 4.315 3.505 4.315 3.505 3.285 2.555 3.285 2.555 3.685 2.325 3.685  ;
        POLYGON 6.105 3.045 8.375 3.045 8.375 3.855 8.145 3.855 8.145 3.275 6.335 3.275 6.335 3.855 6.105 3.855  ;
        POLYGON 5.085 2.765 5.445 2.765 5.445 1.225 5.675 1.225 5.675 2.585 9.59 2.585 9.59 2.815 5.67 2.815 5.67 2.995 5.315 2.995 5.315 3.685 5.085 3.685  ;
        POLYGON 6.67 1.95 9.635 1.95 9.635 1.225 9.865 1.225 9.865 2.13 10.115 2.13 10.115 3.995 9.885 3.995 9.885 2.36 9.64 2.36 9.64 2.18 6.67 2.18  ;
        POLYGON 6.125 1.455 9.175 1.455 9.175 0.765 11.575 0.765 11.575 3.065 11.345 3.065 11.345 0.995 10.55 0.995 10.55 2.025 10.32 2.025 10.32 0.995 9.405 0.995 9.405 1.685 6.355 1.685 6.355 2.025 6.125 2.025  ;
        POLYGON 11.9 1.225 12.155 1.225 12.155 3.525 11.9 3.525  ;
        POLYGON 10.78 1.225 11.01 1.225 11.01 3.185 11.135 3.185 11.135 3.765 14.72 3.765 14.72 2.725 14.95 2.725 14.95 3.995 10.78 3.995  ;
        POLYGON 12.58 2.725 12.81 2.725 12.81 3.295 14.26 3.295 14.26 2.265 15.44 2.265 15.44 1.315 15.67 1.315 15.67 1.975 15.93 1.975 15.93 2.495 14.49 2.495 14.49 3.525 12.58 3.525  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1
