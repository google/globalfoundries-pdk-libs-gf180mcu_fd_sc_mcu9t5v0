* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(((A1 + A2) * (B1 + B2)) * (C1 + C2))
M_i_5 net_1 C2 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4 VSS C1 net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2 net_1 B1 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3 net_0 B2 net_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1 ZN A2 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0 net_0 A1 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_11 net_4 C2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_10 ZN C1 net_4 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8 net_3 B1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9 VDD B2 net_3 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_7 net_2 A2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6 ZN A1 net_2 VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
