* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__invz_4 EN I ZN VDD VNW VPW VSS
*.PININFO EN:I I:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!I
M_mn VSS EN NEN VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn8 NI_N NEN VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn21 NI_P EN NI_N VPW nfet_05v0 W=1.320000U L=0.600000U
M_Mn_inv VSS I NI VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn17 NI_N NI VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn17_9 VSS NI NI_N VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3 ZN NI_N VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_1 VSS NI_N ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_49 ZN NI_N VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_1_25 VSS NI_N ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_mp VDD EN NEN VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp7 NI_P EN VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp22 NI_N NEN NI_P VNW pfet_05v0 W=1.800000U L=0.500000U
M_Mp_inv VDD I NI VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp14 NI_P NI VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp14_10 VDD NI NI_P VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4 ZN NI_P VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_12 VDD NI_P ZN VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_56 ZN NI_P VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_12_57 VDD NI_P ZN VNW pfet_05v0 W=1.800000U L=0.500000U
.ENDS
