# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

##################################################################################
#
#           GLOBALFOUNDRIES
#
##################################################################################
#
# 180MCU Tech LEF File
# based on DRM DM-000013-01 Rev 13
# TFG-Version: 2.1.9
# Date: February 2018
#-------------------------------------------------------
# metal stack option: 3LM_1TM_11K
# Preferred routing directions:
# vertical:   Metal2 
# horizontal: Metal1 Metal3
#------------------------------------------------------
# This Techfile contains not correct Parasitic Information.
# USE Appropriate parasitic files for Parasitic Extraction.
#------------------------------------------------------

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE GF018hv5v_green_sc9
  SYMMETRY X Y ;
  CLASS core ;
  SIZE 0.56 BY 5.04 ;
END GF018hv5v_green_sc9

UNITS
    DATABASE MICRONS 2000  ;
    CAPACITANCE PICOFARADS 1 ;
    CURRENT MILLIAMPS 1 ;
    RESISTANCE OHMS 1 ;
END UNITS

PROPERTYDEFINITIONS
  LAYER LEF58_EOLENCLOSURE STRING ;
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

MANUFACTURINGGRID 0.0050 ;
CLEARANCEMEASURE EUCLIDEAN ;
USEMINSPACING OBS ON ;

LAYER Poly2
    TYPE MASTERSLICE ;
END Poly2

LAYER CON
    TYPE CUT ;
END CON



LAYER Metal1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;

    PITCH 0.56 ;
    OFFSET 0.0 ;  

    MINWIDTH 0.230 ;                   # Mn.1  (n=1)
    WIDTH 0.230 ;                      # Mn.1  (n=1)
    SPACING 0.230  ;                   # Mn.2a (n=1)
    SPACING 0.300 RANGE 10.005 999.00 ; # Mn.2b
    AREA 0.1444 ;                      # Mn.3

    THICKNESS 0.54 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;

    DCCURRENTDENSITY AVERAGE 0.67 ;
    ACCURRENTDENSITY AVERAGE 1.00 ;

    CAPACITANCE CPERSQDIST 0.0000394 ;
    RESISTANCE RPERSQ 0.090000 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END Metal1


LAYER Via1
  TYPE CUT ;
  SPACING 0.26 ;
  WIDTH   0.26 ;

  ENCLOSURE BELOW 0.00 0.06 ;
  ENCLOSURE ABOVE 0.01 0.06 ;
  PROPERTY LEF58_EOLENCLOSURE "
  	EOLENCLOSURE 0.34 0.06 ;" ; 

  ARRAYSPACING CUTSPACING 0.36 ARRAYCUTS 4 SPACING 0.36 ; # Vn.2b

  ACCURRENTDENSITY AVERAGE 0.28 ;
  DCCURRENTDENSITY AVERAGE 0.18 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNAAREARATIO 20.0 ;
END Via1


LAYER Metal2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;

    PITCH 0.56 ;
    OFFSET 0.0 ;  

    MINWIDTH 0.280 ;
    WIDTH 0.280 ;                        # Mn.1  (n>1)
    SPACING 0.280 ;                      # Mn.2a (n>1)
    SPACING 0.300 RANGE 10.005 999.00 ;  # Mn.2b
    AREA 0.1444 ;                        # Mn.3

    THICKNESS 0.54 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO 400 ;
    ANTENNAGATEPLUSDIFF 2 ;

    DCCURRENTDENSITY AVERAGE 0.67 ;
    ACCURRENTDENSITY AVERAGE 1.00 ;

    CAPACITANCE CPERSQDIST 0.0000394 ;
    RESISTANCE RPERSQ 0.090000 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END Metal2


LAYER Via2
  TYPE CUT ;
  SPACING 0.26 ;
  WIDTH   0.26 ;

  ENCLOSURE BELOW 0.01 0.06 ;
  ENCLOSURE ABOVE 0.01 0.06 ;

  # a bit conservative for Vn.3/4a without considering the protrusion length of 0.28
  PROPERTY LEF58_EOLENCLOSURE " EOLENCLOSURE 0.34 0.06 ; " ;

  ARRAYSPACING CUTSPACING 0.36 ARRAYCUTS 4 SPACING 0.36 ; # Vn.2b

  ACCURRENTDENSITY AVERAGE 0.28 ;
  DCCURRENTDENSITY AVERAGE 0.18 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNAAREARATIO 20.0 ;
END Via2



LAYER Metal3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;

    OFFSET 0.0 ;  


    PITCH 0.9 ;
    MINWIDTH 0.440 ;
    WIDTH   0.440 ;                      # MT.1
    AREA    0.5625 ;                     # MT.4
    SPACING 0.460 ;                      # MT.2a
    SPACING 0.600 RANGE 10.005 999.00 ;  # MT.2b

    DCCURRENTDENSITY AVERAGE 1.5 ;
    ACCURRENTDENSITY AVERAGE 2.2 ;
    RESISTANCE RPERSQ 0.04000 ;

    THICKNESS 1.19 ;

    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO 400 ;
    ANTENNAGATEPLUSDIFF 2 ;

    CAPACITANCE CPERSQDIST 0.0000394 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END Metal3



LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER PR_bndry
    TYPE MASTERSLICE ;
END PR_bndry


#------------------------------------------------------------
#  Via1 VIA SECTION 
#------------------------------------------------------------
 VIA Via1_HH  DEFAULT
 LAYER Via1 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal1 ;
 RECT -0.190 -0.130 0.190 0.130 ;
 LAYER Metal2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via1_HH 
 
 VIA Via1_HV  DEFAULT
 LAYER Via1 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal1 ;
 RECT -0.190 -0.130 0.190 0.130 ;
 LAYER Metal2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via1_HV 
 
 VIA Via1_VH  DEFAULT
 LAYER Via1 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal1 ;
 RECT -0.130 -0.190 0.130 0.190 ;
 LAYER Metal2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via1_VH 
 
 VIA Via1_VV  DEFAULT
 LAYER Via1 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal1 ;
 RECT -0.130 -0.190 0.130 0.190 ;
 LAYER Metal2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via1_VV 
 
 VIA Via1_2CUT_H
 LAYER Via1 ;
 RECT -0.390 -0.130 -0.130 0.130 ;
 RECT 0.130 -0.130 0.390 0.130 ;
 LAYER Metal1 ;
 RECT -0.450 -0.130 0.450 0.130 ;
 LAYER Metal2 ;
 RECT -0.400 -0.190 0.400 0.190 ;
 END Via1_2CUT_H
 
 VIA Via1_2CUT_V
 LAYER Via1 ;
 RECT -0.130 -0.390 0.130 -0.130 ;
 RECT -0.130 0.130 0.130 0.390 ;
 LAYER Metal1 ;
 RECT -0.190 -0.390 0.190 0.390 ;
 LAYER Metal2 ;
 RECT -0.140 -0.450 0.140 0.450 ;
 END Via1_2CUT_V
 
 VIA Via1_2X2_0_60_10_60_H_H  DEFAULT
 LAYER Via1 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal1 ;
 RECT -0.450 -0.390 0.450 0.390 ;
 LAYER Metal2 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via1_2X2_0_60_10_60_H_H 
 
 VIA Via1_2X2_0_60_10_60_H_V  DEFAULT
 LAYER Via1 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal1 ;
 RECT -0.450 -0.390 0.450 0.390 ;
 LAYER Metal2 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via1_2X2_0_60_10_60_H_V 
 
 VIA Via1_2X2_0_60_10_60_V_H  DEFAULT
 LAYER Via1 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal1 ;
 RECT -0.390 -0.450 0.390 0.450 ;
 LAYER Metal2 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via1_2X2_0_60_10_60_V_H 
 
 VIA Via1_2X2_0_60_10_60_V_V  DEFAULT
 LAYER Via1 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal1 ;
 RECT -0.390 -0.450 0.390 0.450 ;
 LAYER Metal2 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via1_2X2_0_60_10_60_V_V 
 
VIARULE Via1_GEN_HH GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.060 0.000 ;
  LAYER Metal2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via1 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via1_GEN_HH

VIARULE Via1_GEN_HV GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.060 0.000 ;
  LAYER Metal2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via1 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via1_GEN_HV

VIARULE Via1_GEN_VH GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.000 0.060 ;
  LAYER Metal2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via1 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via1_GEN_VH

VIARULE Via1_GEN_VV GENERATE
  LAYER Metal1 ;
    ENCLOSURE 0.000 0.060 ;
  LAYER Metal2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via1 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via1_GEN_VV

 VIA Via1_4X4H_HH_DEFAULT  DEFAULT
 LAYER Via1 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal1 ;
 RECT -1.120 -1.060 1.120 1.060 ;
 LAYER Metal2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via1_4X4H_HH_DEFAULT 
 
 VIA Via1_4X4H_HV_DEFAULT  DEFAULT
 LAYER Via1 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal1 ;
 RECT -1.120 -1.060 1.120 1.060 ;
 LAYER Metal2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via1_4X4H_HV_DEFAULT 
 
 VIA Via1_4X4H_VH_DEFAULT  DEFAULT
 LAYER Via1 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal1 ;
 RECT -1.060 -1.120 1.060 1.120 ;
 LAYER Metal2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via1_4X4H_VH_DEFAULT 
 
 VIA Via1_4X4H_VV_DEFAULT  DEFAULT
 LAYER Via1 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal1 ;
 RECT -1.060 -1.120 1.060 1.120 ;
 LAYER Metal2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via1_4X4H_VV_DEFAULT 
 
#------------------------------------------------------------
#  Via2 VIA SECTION 
#------------------------------------------------------------
 VIA Via2_HH  DEFAULT
 LAYER Via2 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER Metal3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via2_HH 
 
 VIA Via2_HV  DEFAULT
 LAYER Via2 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER Metal3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via2_HV 
 
 VIA Via2_VH  DEFAULT
 LAYER Via2 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER Metal3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 RESISTANCE 4.500 ;
 END Via2_VH 
 
 VIA Via2_VV  DEFAULT
 LAYER Via2 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER Metal2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER Metal3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 RESISTANCE 4.500 ;
 END Via2_VV 
 
 VIA Via2_2CUT_H
 LAYER Via2 ;
 RECT -0.390 -0.130 -0.130 0.130 ;
 RECT 0.130 -0.130 0.390 0.130 ;
 LAYER Metal2 ;
 RECT -0.400 -0.190 0.400 0.190 ;
 LAYER Metal3 ;
 RECT -0.450 -0.140 0.450 0.140 ;
 END Via2_2CUT_H
 
 VIA Via2_2CUT_V
 LAYER Via2 ;
 RECT -0.130 -0.390 0.130 -0.130 ;
 RECT -0.130 0.130 0.130 0.390 ;
 LAYER Metal2 ;
 RECT -0.140 -0.450 0.140 0.450 ;
 LAYER Metal3 ;
 RECT -0.190 -0.400 0.190 0.400 ;
 END Via2_2CUT_V
 
 VIA Via2_2X2_10_60_10_60_H_H  DEFAULT
 LAYER Via2 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal2 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 LAYER Metal3 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via2_2X2_10_60_10_60_H_H 
 
 VIA Via2_2X2_10_60_10_60_H_V  DEFAULT
 LAYER Via2 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal2 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 LAYER Metal3 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via2_2X2_10_60_10_60_H_V 
 
 VIA Via2_2X2_10_60_10_60_V_H  DEFAULT
 LAYER Via2 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal2 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 LAYER Metal3 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END Via2_2X2_10_60_10_60_V_H 
 
 VIA Via2_2X2_10_60_10_60_V_V  DEFAULT
 LAYER Via2 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER Metal2 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 LAYER Metal3 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END Via2_2X2_10_60_10_60_V_V 
 
VIARULE Via2_GEN_HH GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Metal3 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via2 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via2_GEN_HH

VIARULE Via2_GEN_HV GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Metal3 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via2 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via2_GEN_HV

VIARULE Via2_GEN_VH GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Metal3 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER Via2 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via2_GEN_VH

VIARULE Via2_GEN_VV GENERATE
  LAYER Metal2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Metal3 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER Via2 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END Via2_GEN_VV

 VIA Via2_4X4H_HH_DEFAULT  DEFAULT
 LAYER Via2 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER Metal3 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via2_4X4H_HH_DEFAULT 
 
 VIA Via2_4X4H_HV_DEFAULT  DEFAULT
 LAYER Via2 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER Metal3 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via2_4X4H_HV_DEFAULT 
 
 VIA Via2_4X4H_VH_DEFAULT  DEFAULT
 LAYER Via2 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER Metal3 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END Via2_4X4H_VH_DEFAULT 
 
 VIA Via2_4X4H_VV_DEFAULT  DEFAULT
 LAYER Via2 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER Metal2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER Metal3 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END Via2_4X4H_VV_DEFAULT 
 

END LIBRARY
