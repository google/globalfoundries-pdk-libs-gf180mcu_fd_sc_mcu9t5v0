* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__oai33_4 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(((A1 + A2) + A3) * ((B1 + B2) + B3))
M_i_4_0 VSS B2 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_5_0 net_0 B3 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_5_1 VSS B3 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4_1 net_0 B2 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4_2 VSS B2 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_5_2 net_0 B3 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_5_3 VSS B3 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4_3 net_0 B2 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_0 VSS B1 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_1 net_0 B1 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_2 VSS B1 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_3 net_0 B1 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0 ZN A1 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_1 net_0 A1 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_2 ZN A1 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_3 net_0 A1 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_3 ZN A2 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_3 net_0 A3 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_2 ZN A3 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_2 net_0 A2 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_1 ZN A2 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_1 net_0 A3 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_0 ZN A3 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1_0 net_0 A2 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_10_0 net_4_0 B2 net_3 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_11_0 VDD B3 net_4_0 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_11_1 net_4_1 B3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_10_1 net_3 B2 net_4_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_10_2 net_4_2 B2 net_3 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_11_2 VDD B3 net_4_2 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_11_3 net_4_3 B3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_10_3 net_3_0 B2 net_4_3 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_0 ZN B1 net_3_0 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_1 net_3 B1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_2 ZN B1 net_3 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9_3 net_3 B1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_0 ZN A1 net_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_1 net_1 A1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_2 ZN A1 net_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_3 net_1_0 A1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_7_3 net_2_0 A2 net_1_0 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8_3 VDD A3 net_2_0 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8_2 net_2_1 A3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_7_2 net_1 A2 net_2_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_7_1 net_2_2 A2 net_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8_1 VDD A3 net_2_2 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8_0 net_2_3 A3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_7_0 net_1 A2 net_2_3 VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
