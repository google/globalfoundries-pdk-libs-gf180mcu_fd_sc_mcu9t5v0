# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyb_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyb_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.64 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.9 0.97 1.9 0.97 2.71 0.71 2.71  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.825 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.74 3.42 8.175 3.42 8.93 3.42 8.93 1.59 6.69 1.59 6.69 0.68 6.92 0.68 6.92 1.21 8.93 1.21 8.93 0.68 9.16 0.68 9.16 4.36 8.93 4.36 8.93 3.65 8.175 3.65 6.97 3.65 6.97 4.36 6.74 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.32 4.59 1.32 4.06 1.55 4.06 1.55 4.59 4.44 4.59 4.79 4.59 4.79 4.06 5.02 4.06 5.02 4.59 7.76 4.59 7.76 3.88 7.99 3.88 7.99 4.59 8.175 4.59 9.95 4.59 9.95 3.88 10.18 3.88 10.18 4.59 10.64 4.59 10.64 5.49 8.175 5.49 4.44 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 10.64 -0.45 10.64 0.45 10.28 0.45 10.28 1.435 10.05 1.435 10.05 0.45 8.04 0.45 8.04 0.965 7.81 0.965 7.81 0.45 5.12 0.45 5.12 0.695 4.89 0.695 4.89 0.45 1.65 0.45 1.65 0.965 1.42 0.965 1.42 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.475 2.94 1.275 2.94 1.275 2.425 2.05 2.425 2.05 1.9 2.335 1.9 2.335 2.655 1.505 2.655 1.505 3.17 0.585 3.17 0.585 4.345 0.245 4.345 0.245 0.68 0.585 0.68 0.585 0.91 0.475 0.91  ;
        POLYGON 1.555 3.395 2.565 3.395 2.565 1.63 1.555 1.63 1.555 1.4 4.44 1.4 4.44 2.71 4.21 2.71 4.21 1.63 2.795 1.63 2.795 3.625 1.555 3.625  ;
        POLYGON 4.79 1.075 5.12 1.075 5.12 2.19 8.175 2.19 8.175 2.42 5.02 2.42 5.02 3.68 4.79 3.68  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyb_4
