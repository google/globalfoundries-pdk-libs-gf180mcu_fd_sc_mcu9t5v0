# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 34.72 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 17.07 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.685 2.215 9.845 2.215 9.845 2.65 0.685 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 18.21 ;
    PORT
      LAYER METAL1 ;
        POLYGON 12.565 2.885 21.1 2.885 22.285 2.885 22.285 2.03 12.565 2.03 12.565 0.68 12.825 0.68 12.825 1.72 14.805 1.72 14.805 0.68 15.035 0.68 15.035 1.72 17.045 1.72 17.045 0.68 17.275 0.68 17.275 1.72 19.285 1.72 19.285 0.68 19.515 0.68 19.515 1.72 21.525 1.72 21.525 0.68 21.755 0.68 21.755 1.72 23.765 1.72 23.765 0.68 23.995 0.68 23.995 1.72 26.005 1.72 26.005 0.68 26.235 0.68 26.235 1.72 28.245 1.72 28.245 0.68 28.475 0.68 28.475 1.72 30.485 1.72 30.485 0.68 30.715 0.68 30.715 1.72 32.725 1.72 32.725 0.68 32.955 0.68 32.955 1.98 23.035 1.98 23.035 2.88 32.425 2.88 32.855 2.88 32.855 4.36 32.625 4.36 32.625 3.32 32.425 3.32 30.615 3.32 30.615 4.36 30.385 4.36 30.385 3.32 28.375 3.32 28.375 4.36 28.145 4.36 28.145 3.32 26.135 3.32 26.135 4.36 25.905 4.36 25.905 3.32 23.895 3.32 23.895 4.36 23.665 4.36 23.665 3.32 21.655 3.32 21.655 4.36 21.425 4.36 21.425 3.32 21.1 3.32 19.415 3.32 19.415 4.36 19.185 4.36 19.185 3.32 17.175 3.32 17.175 4.36 16.945 4.36 16.945 3.32 14.935 3.32 14.935 4.36 14.705 4.36 14.705 3.32 12.795 3.32 12.795 4.36 12.565 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.875 11.575 3.875 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 15.825 4.59 15.825 3.55 16.055 3.55 16.055 4.59 18.065 4.59 18.065 3.55 18.295 3.55 18.295 4.59 20.305 4.59 20.305 3.55 20.535 3.55 20.535 4.59 21.1 4.59 22.545 4.59 22.545 3.55 22.775 3.55 22.775 4.59 24.785 4.59 24.785 3.55 25.015 3.55 25.015 4.59 27.025 4.59 27.025 3.55 27.255 3.55 27.255 4.59 29.265 4.59 29.265 3.55 29.495 3.55 29.495 4.59 31.505 4.59 31.505 3.55 31.735 3.55 31.735 4.59 32.425 4.59 33.745 4.59 33.745 3.55 33.975 3.55 33.975 4.59 34.72 4.59 34.72 5.49 32.425 5.49 21.1 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 34.72 -0.45 34.72 0.45 34.075 0.45 34.075 1.49 33.845 1.49 33.845 0.45 31.835 0.45 31.835 1.49 31.605 1.49 31.605 0.45 29.595 0.45 29.595 1.49 29.365 1.49 29.365 0.45 27.355 0.45 27.355 1.49 27.125 1.49 27.125 0.45 25.115 0.45 25.115 1.49 24.885 1.49 24.885 0.45 22.875 0.45 22.875 1.49 22.645 1.49 22.645 0.45 20.635 0.45 20.635 1.49 20.405 1.49 20.405 0.45 18.395 0.45 18.395 1.49 18.165 1.49 18.165 0.45 16.155 0.45 16.155 1.49 15.925 1.49 15.925 0.45 13.915 0.45 13.915 1.49 13.685 1.49 13.685 0.45 11.675 0.45 11.675 1.49 11.445 1.49 11.445 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.365 2.9 10.225 2.9 10.225 1.975 1.365 1.975 1.365 0.68 1.595 0.68 1.595 1.72 3.605 1.72 3.605 0.68 3.835 0.68 3.835 1.72 5.845 1.72 5.845 0.68 6.075 0.68 6.075 1.72 8.085 1.72 8.085 0.68 8.315 0.68 8.315 1.72 10.325 1.72 10.325 0.68 10.555 0.68 10.555 2.27 21.1 2.27 21.1 2.65 10.555 2.65 10.555 4.36 10.225 4.36 10.225 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
        POLYGON 23.265 2.215 32.425 2.215 32.425 2.65 23.265 2.65  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_20
