# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.698 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.87 2.33 2.09 2.33 2.09 2.71 0.87 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.849 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.63 1.745 4.99 1.745 4.99 2.15 4.63 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.64 0.84 7.13 0.84 7.13 1.65 6.87 1.65 6.87 3.685 6.64 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.635 1.595 3.635 1.595 4.59 5.44 4.59 5.44 3.875 5.67 3.875 5.67 4.59 6.345 4.59 6.385 4.59 7.28 4.59 7.28 5.49 6.385 5.49 6.345 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 5.89 0.45 5.89 0.69 5.66 0.69 5.66 0.45 1.595 0.45 1.595 1.425 1.365 1.425 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 1.315 0.475 1.315 0.475 1.83 2.86 1.83 2.86 2.815 2.895 2.815 2.895 3.155 2.63 3.155 2.63 2.06 0.575 2.06 0.575 4.285 0.245 4.285  ;
        POLYGON 2.385 3.475 2.615 3.475 2.615 4.055 4.17 4.055 4.17 1.6 3.55 1.6 3.55 1.37 4.4 1.37 4.4 2.47 6.345 2.47 6.345 2.7 4.65 2.7 4.65 4.285 2.385 4.285  ;
        POLYGON 2.485 0.72 5.43 0.72 5.43 0.92 6.385 0.92 6.385 2.055 5.305 2.055 5.305 1.115 3.32 1.115 3.32 1.83 3.635 1.83 3.635 3.815 3.405 3.815 3.405 2.06 3.09 2.06 3.09 0.95 2.715 0.95 2.715 1.425 2.485 1.425  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_1
