# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 11.76 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.63 3.39 2.63 3.62 2.63 3.62 2.17 4.51 2.17 4.51 2.4 3.85 2.4 3.85 2.86 3.39 2.86 1.83 2.86  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.985 1.77 0.985 3.09 3.39 3.09 4.625 3.09 4.625 2.6 5.245 2.6 5.245 2.115 5.475 2.115 5.475 2.83 4.855 2.83 4.855 3.32 3.39 3.32 0.755 3.32 0.755 2.455 0.71 2.455  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 2.89 7.665 2.89 7.665 0.68 7.895 0.68 7.895 1.72 9.905 1.72 9.905 0.68 10.135 0.68 10.135 3.685 9.855 3.685 9.855 1.95 7.895 1.95 7.895 3.685 7.665 3.685 7.665 3.27 7.43 3.27  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.665 4.59 2.665 3.875 2.895 3.875 2.895 4.59 3.39 4.59 6.11 4.59 6.645 4.59 6.645 3.875 6.875 3.875 6.875 4.59 7.315 4.59 8.735 4.59 8.735 3.875 8.965 3.875 8.965 4.59 10.925 4.59 10.925 2.875 11.155 2.875 11.155 4.59 11.76 4.59 11.76 5.49 7.315 5.49 6.11 5.49 3.39 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 11.76 -0.45 11.76 0.45 11.255 0.45 11.255 1.49 11.025 1.49 11.025 0.45 9.015 0.45 9.015 1.49 8.785 1.49 8.785 0.45 6.775 0.45 6.775 1.425 6.545 1.425 6.545 0.45 6.055 0.45 6.055 1.425 5.825 1.425 5.825 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.02 0.245 1.02 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.25 1.31 1.365 1.31 1.365 0.68 1.595 0.68 1.595 1.31 2.55 1.31 2.55 2.17 3.39 2.17 3.39 2.4 2.32 2.4 2.32 1.54 0.48 1.54 0.48 2.875 0.525 2.875 0.525 3.215 0.25 3.215  ;
        POLYGON 3.785 3.55 4.015 3.55 4.015 4.13 6.11 4.13 6.11 4.36 3.785 4.36  ;
        POLYGON 4.75 3.55 5.705 3.55 5.705 1.885 3.785 1.885 3.785 0.68 4.015 0.68 4.015 1.655 7.315 1.655 7.315 2.455 7.085 2.455 7.085 1.885 5.935 1.885 5.935 3.78 4.75 3.78  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor2_4
