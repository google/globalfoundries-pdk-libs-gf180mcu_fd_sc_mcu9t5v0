# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nor4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.465 2.215 17.46 2.215 17.46 2.71 13.465 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.87 1.755 20.01 1.755 20.01 2.555 19.55 2.555 19.55 1.985 11.1 1.985 11.1 2.555 10.87 2.555  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.33 1.77 1.33 2.785 4.59 2.785 4.59 2.215 4.82 2.215 4.82 2.785 7.47 2.785 7.47 2.27 9.715 2.27 9.715 2.5 7.7 2.5 7.7 3.015 1.1 3.015 1.1 2.15 0.71 2.15  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.48 1.755 7.24 1.755 7.24 2.555 6.78 2.555 6.78 1.985 3.71 1.985 3.71 2.555 3.48 2.555  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.3894 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.89 3.09 20.405 3.09 20.405 1.59 20.175 1.59 20.175 1.455 6.52 1.455 6.52 0.91 5.91 0.91 5.91 1.455 1.68 1.455 1.68 0.68 1.91 0.68 1.91 1.225 3.92 1.225 3.92 0.68 4.15 0.68 4.15 1.225 5.68 1.225 5.68 0.68 6.75 0.68 6.75 1.225 8.76 1.225 8.76 0.68 8.99 0.68 8.99 1.225 11.36 1.225 11.36 0.68 11.59 0.68 11.59 1.225 13.96 1.225 13.96 0.68 14.19 0.68 14.19 1.225 16.56 1.225 16.56 0.68 16.79 0.68 16.79 1.225 19.16 1.225 19.16 0.68 19.39 0.68 19.39 1.21 20.635 1.21 20.635 3.32 18.04 3.32 18.04 3.9 17.81 3.9 17.81 3.32 13.12 3.32 13.12 3.9 12.89 3.9  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.75 4.59 2.75 3.705 2.98 3.705 2.98 4.59 7.59 4.59 7.59 3.705 7.82 3.705 7.82 4.59 20.59 4.59 21.28 4.59 21.28 5.49 20.59 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.69 0.45 20.69 0.98 20.46 0.98 20.46 0.45 18.09 0.45 18.09 0.995 17.86 0.995 17.86 0.45 15.49 0.45 15.49 0.97 15.26 0.97 15.26 0.45 12.89 0.45 12.89 0.995 12.66 0.995 12.66 0.45 10.29 0.45 10.29 0.995 10.06 0.995 10.06 0.45 7.87 0.45 7.87 0.995 7.64 0.995 7.64 0.45 5.45 0.45 5.45 0.995 5.22 0.995 5.22 0.45 3.03 0.45 3.03 0.995 2.8 0.995 2.8 0.45 0.79 0.45 0.79 0.995 0.56 0.995 0.56 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.66 3.55 0.89 3.55 0.89 4.13 2.29 4.13 2.29 3.245 8.28 3.245 8.28 4.13 15.21 4.13 15.21 3.55 15.44 3.55 15.44 4.13 20.36 4.13 20.36 3.55 20.59 3.55 20.59 4.36 8.05 4.36 8.05 3.475 5.4 3.475 5.4 4.36 5.17 4.36 5.17 3.475 2.52 3.475 2.52 4.36 0.66 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nor4_4
