# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.04 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER METAL1 ;
        POLYGON 16.95 1.21 17.21 1.21 17.21 2.03 16.95 2.03  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER METAL1 ;
        POLYGON 13.59 1.77 13.85 1.77 13.85 2.39 13.59 2.39  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.05 1.015 2.05 1.015 3.27 0.71 3.27  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.625 2.05 4.89 2.05 4.89 2.71 4.625 2.71  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.36 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.285 1.77 3.815 1.77 3.815 2.26 3.51 2.26 3.51 2 2.515 2 2.515 2.39 2.285 2.39  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.24 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.56 1.69 9.79 1.69 9.79 1.77 10.23 1.77 10.83 1.77 10.83 2.83 10.6 2.83 10.6 2.15 10.23 2.15 9.56 2.15  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0816 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.31 1.2 6.755 1.2 6.755 3.38 6.31 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.25 4.59 0.25 3.08 0.48 3.08 0.48 4.59 1.595 4.59 5.285 4.59 5.285 4.07 5.515 4.07 5.515 4.59 7.545 4.59 7.545 3.08 7.775 3.08 7.775 4.59 9.005 4.59 10.23 4.59 13 4.59 13 3.08 13.23 3.08 13.23 4.59 15.43 4.59 17.34 4.59 17.34 3.08 17.57 3.08 17.57 4.59 18.79 4.59 19.04 4.59 19.04 5.49 18.79 5.49 15.43 5.49 10.23 5.49 9.005 5.49 1.595 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 19.04 -0.45 19.04 0.45 17.67 0.45 17.67 1.54 17.44 1.54 17.44 0.45 13.19 0.45 13.19 1.54 12.96 1.54 12.96 0.45 7.875 0.45 7.875 1.54 7.645 1.54 7.645 0.45 5.635 0.45 5.635 1.54 5.405 1.54 5.405 0.45 0.475 0.45 0.475 1.54 0.245 1.54 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.365 1.2 1.595 1.2 1.595 3.89 1.365 3.89  ;
        POLYGON 4.045 1.615 4.285 1.615 4.285 1.2 4.515 1.2 4.515 1.845 4.275 1.845 4.275 3.38 4.045 3.38  ;
        POLYGON 2.055 3.61 2.725 3.61 2.725 3.08 2.955 3.08 2.955 3.61 7.085 3.61 7.085 2.62 8.64 2.62 8.64 1.21 8.87 1.21 8.87 3.08 9.005 3.08 9.005 3.89 8.64 3.89 8.64 2.85 7.315 2.85 7.315 3.84 2.955 3.84 2.955 3.89 1.825 3.89 1.825 1.255 3.45 1.255 3.45 1.485 2.055 1.485  ;
        POLYGON 7.105 1.77 8.18 1.77 8.18 0.75 10.23 0.75 10.23 1.54 10 1.54 10 0.98 9.33 0.98 9.33 2.36 9.465 2.36 9.465 3.66 9.95 3.66 9.95 3.08 10.18 3.08 10.18 3.89 9.235 3.89 9.235 2.57 9.1 2.57 9.1 0.98 8.41 0.98 8.41 2 7.335 2 7.335 2.39 7.105 2.39  ;
        POLYGON 11.68 1.2 12.21 1.2 12.21 3.89 11.68 3.89  ;
        POLYGON 14.08 1.2 14.31 1.2 14.31 3.89 14.08 3.89  ;
        POLYGON 11.12 1.2 11.41 1.2 11.41 4.12 12.54 4.12 12.54 2.62 13.69 2.62 13.69 4.12 15.17 4.12 15.17 1.2 15.43 1.2 15.43 4.35 13.46 4.35 13.46 2.85 12.77 2.85 12.77 4.35 11.12 4.35  ;
        POLYGON 15.7 1.255 16.605 1.255 16.605 1.485 15.93 1.485 15.93 2.665 16.42 2.665 16.42 3.89 16.19 3.89 16.19 2.895 15.7 2.895  ;
        POLYGON 16.16 2.05 16.72 2.05 16.72 2.26 18.56 2.26 18.56 1.2 18.79 1.2 18.79 3.89 18.46 3.89 18.46 2.49 16.57 2.49 16.57 2.435 16.16 2.435  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_2
