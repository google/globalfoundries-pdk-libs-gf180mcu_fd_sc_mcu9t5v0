* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(A1 + A2)
M_i_1_3 ZN A2 VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_0_3 VSS A1 ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_0_2 ZN A1 VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_1_2 VSS A2 ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_1_1 ZN A2 VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_0_1 VSS A1 ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_0_0 ZN A1 VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_1_0 VSS A2 ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_3_3 net_0_0 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_2_3 ZN A1 net_0_0 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_2_2 net_0_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 VDD A2 net_0_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 net_0_2 A2 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_2_1 ZN A1 net_0_2 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_2_0 net_0_3 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 VDD A2 net_0_3 VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
