# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 3.92 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.21 3.21 1.21 3.21 2.15 2.95 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.71 1.83 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.33 1.105 2.33 1.105 3.27 0.71 3.27  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9824 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 3.55 2.95 3.55 2.95 2.89 3.44 2.89 3.44 0.845 3.67 0.845 3.67 3.83 1.63 3.83 1.63 4.36 1.4 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.38 4.59 0.38 3.59 0.61 3.59 0.61 4.59 2.42 4.59 2.42 4.06 2.65 4.06 2.65 4.59 3.92 4.59 3.92 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 3.92 -0.45 3.92 0.45 0.61 0.45 0.61 1.165 0.38 1.165 0.38 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand3_1
