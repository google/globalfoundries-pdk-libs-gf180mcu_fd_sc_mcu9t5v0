# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__latrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.36 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.5 1.77 3.5 2.195 3.21 2.195 3.21 2.71 2.95 2.71  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.97 1.965 1.83 1.965 1.83 1.31 4.285 1.31 4.285 1.89 4.755 1.89 4.755 2.875 5.37 2.875 5.37 3.105 4.525 3.105 4.525 2.12 4.055 2.12 4.055 1.54 2.09 1.54 2.09 2.71 1.83 2.71 1.83 2.195 0.97 2.195  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.34 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.375 1.77 2.65 1.77 2.65 2.71 2.375 2.71  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.55 1.77 8.985 1.77 8.985 2.71 8.55 2.71  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.265 3.42 13.515 3.42 13.515 0.845 13.745 0.845 13.745 1.92 15.27 1.92 15.27 1.21 15.755 1.21 15.755 0.845 15.985 0.845 15.985 1.655 15.53 1.655 15.53 2.15 13.745 2.15 13.745 3.42 15.535 3.42 15.535 4.29 15.305 4.29 15.305 3.65 13.495 3.65 13.495 4.29 13.265 4.29  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.305 4.59 1.305 3.48 1.535 3.48 1.535 4.59 3.045 4.59 3.045 4.12 3.275 4.12 3.275 4.59 6.565 4.59 6.565 3.48 6.795 3.48 6.795 4.59 7.535 4.59 8.785 4.59 8.785 3.65 9.015 3.65 9.015 4.59 10.205 4.59 10.205 3.88 10.435 3.88 10.435 4.59 11.065 4.59 12.245 4.59 12.245 3.88 12.475 3.88 12.475 4.59 12.915 4.59 14.285 4.59 14.285 3.88 14.515 3.88 14.515 4.59 16.325 4.59 16.325 3.88 16.555 3.88 16.555 4.59 17.36 4.59 17.36 5.49 12.915 5.49 11.065 5.49 7.535 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.36 -0.45 17.36 0.45 17.105 0.45 17.105 1.165 16.875 1.165 16.875 0.45 14.865 0.45 14.865 1.165 14.635 1.165 14.635 0.45 12.625 0.45 12.625 1.165 12.395 1.165 12.395 0.45 10.385 0.45 10.385 1.165 10.155 1.165 10.155 0.45 7.58 0.45 7.58 1.08 7.24 1.08 7.24 0.45 1.8 0.45 1.8 1.08 1.46 1.08 1.46 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.285 0.795 0.625 0.795 0.625 2.94 4.065 2.94 4.065 2.38 4.295 2.38 4.295 3.17 0.515 3.17 0.515 4.29 0.285 4.29  ;
        POLYGON 2.025 3.48 4.82 3.48 4.82 3.335 5.6 3.335 5.6 2.655 5.535 2.655 5.535 1.135 4.495 1.135 4.495 0.795 5.765 0.795 5.765 2.49 7.305 2.49 7.305 1.935 7.535 1.935 7.535 2.72 5.83 2.72 5.83 3.565 5.035 3.565 5.035 4.29 4.805 4.29 4.805 3.71 2.255 3.71 2.255 4.29 2.025 4.29  ;
        POLYGON 7.765 3.19 9.435 3.19 9.435 1.54 6.365 1.54 6.365 2.26 6.135 2.26 6.135 1.31 9.435 1.31 9.435 0.795 9.665 0.795 9.665 1.91 11.065 1.91 11.065 2.25 9.665 2.25 9.665 3.42 7.995 3.42 7.995 4.29 7.765 4.29  ;
        POLYGON 11.225 2.53 12.685 2.53 12.685 1.655 11.275 1.655 11.275 0.845 11.505 0.845 11.505 1.425 12.915 1.425 12.915 2.76 11.455 2.76 11.455 4.29 11.225 4.29  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrsnq_4
