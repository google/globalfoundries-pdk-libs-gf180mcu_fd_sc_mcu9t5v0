# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nand3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.865 1.21 3.21 1.21 3.21 2.15 2.865 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.79 2.38 4.63 2.38 4.63 1.21 4.995 1.21 4.995 2.61 1.79 2.61  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.77 1.92 1.27 1.92 1.27 1.915 1.53 1.915 1.53 2.84 5.74 2.84 5.74 2.07 6.015 2.07 6.015 3.07 1.3 3.07 1.3 2.15 0.77 2.15  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.964 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.41 3.3 5.575 3.3 5.575 4.11 5.345 4.11 5.345 3.53 3.535 3.53 3.535 4.11 3.305 4.11 3.305 3.53 1.495 3.53 1.495 4.11 1.265 4.11 1.265 3.53 0.15 3.53 0.15 0.865 0.87 0.865 0.87 0.75 3.59 0.75 3.59 0.98 1.07 0.98 1.07 1.095 0.41 1.095  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 4.23 0.475 4.23 0.475 4.59 2.285 4.59 2.285 3.76 2.515 3.76 2.515 4.59 4.325 4.59 4.325 3.76 4.555 3.76 4.555 4.59 6.365 4.59 6.365 3.76 6.595 3.76 6.595 4.59 7.28 4.59 7.28 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 6.595 0.45 6.595 1.16 6.365 1.16 6.365 0.45 0.67 0.45 0.67 0.635 0.33 0.635 0.33 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand3_2
