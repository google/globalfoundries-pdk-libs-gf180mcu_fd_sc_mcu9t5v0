# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyd_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyd_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 16.24 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.77 0.99 1.77 0.99 2.57 0.65 2.57  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.821 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.53 4.07 14.535 4.07 14.535 3.135 15.125 3.135 15.355 3.135 15.355 1.82 14.635 1.82 14.635 0.845 14.865 0.845 14.865 1.59 15.585 1.59 15.585 3.365 15.125 3.365 14.765 3.365 14.765 4.36 13.53 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.925 1.495 3.925 1.495 4.59 4.385 4.59 4.735 4.59 4.735 3.925 4.965 3.925 4.965 4.59 8.385 4.59 8.735 4.59 8.735 3.925 8.965 3.925 8.965 4.59 12.385 4.59 12.735 4.59 12.735 3.925 12.965 3.925 12.965 4.59 15.125 4.59 15.655 4.59 15.655 3.585 15.885 3.585 15.885 4.59 16.24 4.59 16.24 5.49 15.125 5.49 12.385 5.49 8.385 5.49 4.385 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 16.24 -0.45 16.24 0.45 15.985 0.45 15.985 1.435 15.755 1.435 15.755 0.45 13.065 0.45 13.065 0.695 12.835 0.695 12.835 0.45 9.065 0.45 9.065 0.92 8.835 0.92 8.835 0.45 5.065 0.45 5.065 0.69 4.835 0.69 4.835 0.45 1.595 0.45 1.595 0.965 1.365 0.965 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.8 1.995 2.8 1.995 2.22 2.225 2.22 2.225 3.03 0.475 3.03 0.475 4.265 0.19 4.265 0.19 0.68 0.53 0.68 0.53 0.91 0.42 0.91  ;
        POLYGON 1.5 3.26 4.155 3.26 4.155 1.63 1.5 1.63 1.5 1.4 4.385 1.4 4.385 3.49 1.5 3.49  ;
        POLYGON 4.735 1.07 5.065 1.07 5.065 1.815 6.225 1.815 6.225 2.625 4.965 2.625 4.965 3.545 4.735 3.545  ;
        POLYGON 5.555 2.855 8.155 2.855 8.155 1.585 5.555 1.585 5.555 1.07 5.785 1.07 5.785 1.355 8.385 1.355 8.385 3.085 5.785 3.085 5.785 3.545 5.555 3.545  ;
        POLYGON 8.735 1.3 9.065 1.3 9.065 1.815 10.225 1.815 10.225 2.625 8.965 2.625 8.965 3.545 8.735 3.545  ;
        POLYGON 9.555 2.855 12.155 2.855 12.155 1.585 9.5 1.585 9.5 1.355 12.385 1.355 12.385 3.085 9.785 3.085 9.785 3.545 9.555 3.545  ;
        POLYGON 12.735 1.075 13.065 1.075 13.065 2.05 15.125 2.05 15.125 2.39 12.965 2.39 12.965 3.545 12.735 3.545  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyd_2
