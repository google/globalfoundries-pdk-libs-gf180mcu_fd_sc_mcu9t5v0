# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 22.96 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 2.33 4.33 2.33 4.33 2.71 3.51 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.63 1.77 18.89 1.77 18.89 2.71 18.63 2.71  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 2.33 0.97 2.33 0.97 2.71 0.15 2.71  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 2.33 2.09 2.33 2.09 2.71 1.27 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 2.33 7.13 2.33 7.13 2.71 6.31 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.87 0.845 21.33 0.845 21.33 4.25 20.87 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 3.44 1.545 3.44 1.545 4.59 5.085 4.59 5.085 3.44 5.315 3.44 5.315 4.59 7.18 4.59 7.18 4.03 7.52 4.03 7.52 4.59 9.38 4.59 9.82 4.59 12.155 4.59 12.155 3.91 12.385 3.91 12.385 4.59 13.405 4.59 13.955 4.59 13.955 3.44 14.185 3.44 14.185 4.59 14.31 4.59 15.205 4.59 18.2 4.59 18.2 3.91 18.43 3.91 18.43 4.59 19.91 4.59 20.24 4.59 20.24 3.44 20.47 3.44 20.47 4.59 20.63 4.59 22.12 4.59 22.12 3.44 22.35 3.44 22.35 4.59 22.96 4.59 22.96 5.49 20.63 5.49 19.91 5.49 15.205 5.49 14.31 5.49 13.405 5.49 9.82 5.49 9.38 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 22.96 -0.45 22.96 0.45 22.4 0.45 22.4 1.655 22.17 1.655 22.17 0.45 18.43 0.45 18.43 1.275 18.2 1.275 18.2 0.45 13.495 0.45 13.495 1.44 13.265 1.44 13.265 0.45 7.515 0.45 7.515 1.18 7.285 1.18 7.285 0.45 5.68 0.45 5.68 0.53 5.45 0.53 5.45 0.45 1.595 0.45 1.595 1.285 1.365 1.285 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.295 2.98 2.545 2.98 2.545 2.1 0.245 2.1 0.245 0.945 0.475 0.945 0.475 1.87 4.835 1.87 4.835 2.635 4.605 2.635 4.605 2.1 2.775 2.1 2.775 3.21 0.525 3.21 0.525 4.25 0.295 4.25  ;
        POLYGON 6.16 3.01 7.725 3.01 7.725 2.1 6.165 2.1 6.165 1.21 6.395 1.21 6.395 1.87 7.955 1.87 7.955 3.24 6.16 3.24  ;
        POLYGON 3.325 0.76 6.025 0.76 6.025 0.75 6.855 0.75 6.855 1.41 7.945 1.41 7.945 0.68 9.355 0.68 9.355 1.275 9.125 1.275 9.125 0.91 8.175 0.91 8.175 1.64 6.625 1.64 6.625 0.98 6.095 0.98 6.095 0.99 3.555 0.99 3.555 1.285 3.325 1.285  ;
        POLYGON 3.325 2.98 5.775 2.98 5.775 3.525 9.38 3.525 9.38 3.755 5.545 3.755 5.545 3.21 3.555 3.21 3.555 4.25 3.325 4.25  ;
        POLYGON 8.305 2.39 8.405 2.39 8.405 1.14 8.635 1.14 8.635 2.35 9.82 2.35 9.82 2.58 8.535 2.58 8.535 3.295 8.305 3.295  ;
        POLYGON 11.135 3.44 13.405 3.44 13.405 4.25 13.175 4.25 13.175 3.67 11.365 3.67 11.365 4.25 11.135 4.25  ;
        POLYGON 10.115 0.945 10.475 0.945 10.475 2.865 13.97 2.865 13.97 2.59 14.31 2.59 14.31 3.095 10.345 3.095 10.345 4.25 10.115 4.25  ;
        POLYGON 11.765 2.13 14.605 2.13 14.605 1.155 14.835 1.155 14.835 2.205 15.205 2.205 15.205 4.25 14.975 4.25 14.975 2.435 14.665 2.435 14.665 2.36 11.995 2.36 11.995 2.635 11.765 2.635  ;
        POLYGON 10.825 1.67 14.145 1.67 14.145 0.695 16.83 0.695 16.83 3.15 16.6 3.15 16.6 0.925 15.295 0.925 15.295 1.955 15.065 1.955 15.065 0.925 14.375 0.925 14.375 1.9 11.055 1.9 11.055 2.635 10.825 2.635  ;
        POLYGON 17.08 1.155 17.41 1.155 17.41 3.78 17.08 3.78  ;
        POLYGON 15.67 1.21 16.225 1.21 16.225 4.02 17.74 4.02 17.74 3.45 18.89 3.45 18.89 4.01 19.68 4.01 19.68 2.295 19.91 2.295 19.91 4.24 18.66 4.24 18.66 3.68 17.97 3.68 17.97 4.25 15.995 4.25 15.995 1.44 15.67 1.44  ;
        POLYGON 17.76 2.295 17.99 2.295 17.99 2.94 19.22 2.94 19.22 1.835 20.24 1.835 20.24 0.945 20.63 0.945 20.63 2.635 20.4 2.635 20.4 2.065 19.45 2.065 19.45 3.78 19.22 3.78 19.22 3.17 17.76 3.17  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1
