# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 28.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.19 1.77 27.395 1.77 27.395 2.555 27.165 2.555 27.165 2 22.915 2 22.915 2.145 22.685 2.145 22.685 2 19.66 2 19.66 2.5 19.19 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.7 2.27 22.04 2.27 22.04 2.48 23.11 2.48 23.11 2.27 25.26 2.27 25.26 2.71 21.7 2.71  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.605 2.215 10.835 2.215 10.835 2.89 13.72 2.89 13.72 2.27 14.06 2.27 14.06 3.04 17.995 3.04 18.2 3.04 18.2 2.27 18.54 2.27 18.54 3.27 17.995 3.27 10.605 3.27  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.74 2.27 13.03 2.27 13.03 1.77 14.52 1.77 14.52 2.27 16.25 2.27 16.25 2.5 14.29 2.5 14.29 2 13.29 2 13.29 2.5 12.74 2.5  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.875 2.215 1.105 2.215 1.105 2.785 4.04 2.785 4.04 2.27 4.38 2.27 4.38 2.785 6.85 2.785 6.85 2.27 8.86 2.27 8.86 2.5 7.08 2.5 7.08 3.015 0.875 3.015  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.165 2.215 3.51 2.215 3.51 1.77 4.84 1.77 4.84 2.27 6.62 2.27 6.62 2.5 4.61 2.5 4.61 2 3.77 2 3.77 2.555 3.165 2.555  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 11.5296 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.295 3.245 9.38 3.245 9.38 3.5 17.995 3.5 18.835 3.5 18.835 3.09 27.745 3.09 27.745 1.515 20.005 1.515 20.005 1.14 20.235 1.14 20.235 1.285 22.19 1.285 22.19 1.14 22.53 1.14 22.53 1.285 24.43 1.285 24.43 1.14 24.77 1.14 24.77 1.285 26.67 1.285 26.67 1.14 27.01 1.14 27.01 1.285 27.975 1.285 27.975 4.36 27.745 4.36 27.745 3.32 23.495 3.32 23.495 4.36 23.265 4.36 23.265 3.32 19.065 3.32 19.065 4.36 18.835 4.36 18.835 3.73 17.995 3.73 14.585 3.73 14.585 4.36 12.97 4.36 12.97 3.73 9.385 3.73 9.385 4.36 9.155 4.36 9.155 3.55 4.905 3.55 4.905 4.36 4.675 4.36 4.675 3.475 0.525 3.475 0.525 4.36 0.295 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.705 2.665 3.705 2.665 4.59 6.915 4.59 6.915 3.78 7.145 3.78 7.145 4.59 12.115 4.59 12.115 3.96 12.345 3.96 12.345 4.59 16.595 4.59 16.595 3.96 16.825 3.96 16.825 4.59 17.995 4.59 21.075 4.59 21.075 3.55 21.305 3.55 21.305 4.59 25.555 4.59 25.555 3.55 25.785 3.55 25.785 4.59 28.075 4.59 28.56 4.59 28.56 5.49 28.075 5.49 17.995 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 28.56 -0.45 28.56 0.45 9.435 0.45 9.435 1.525 9.205 1.525 9.205 0.45 7.195 0.45 7.195 1.525 6.965 1.525 6.965 0.45 4.955 0.45 4.955 1.055 4.725 1.055 4.725 0.45 2.715 0.45 2.715 1.525 2.485 1.525 2.485 0.45 0.475 0.45 0.475 1.525 0.245 1.525 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 0.715 1.595 0.715 1.595 1.755 3.05 1.755 3.05 1.295 3.605 1.295 3.605 0.715 3.835 0.715 3.835 1.295 5.845 1.295 5.845 0.715 6.075 0.715 6.075 1.755 8.085 1.755 8.085 0.715 8.315 0.715 8.315 1.755 10.99 1.755 10.99 1.14 11.275 1.14 11.275 1.29 13.23 1.29 13.23 1.14 13.57 1.14 13.57 1.29 15.525 1.29 15.525 1.14 15.81 1.14 15.81 1.755 17.765 1.755 17.765 1.14 17.995 1.14 17.995 1.985 15.58 1.985 15.58 1.52 11.22 1.52 11.22 1.985 5.845 1.985 5.845 1.525 3.28 1.525 3.28 1.985 1.365 1.985  ;
        POLYGON 9.925 0.68 28.075 0.68 28.075 1.055 27.845 1.055 27.845 0.91 25.89 0.91 25.89 1 25.55 1 25.55 0.91 23.65 0.91 23.65 1 23.31 1 23.31 0.91 21.41 0.91 21.41 1 21.07 1 21.07 0.91 19.115 0.91 19.115 1.525 18.885 1.525 18.885 0.91 16.875 0.91 16.875 1.525 16.645 1.525 16.645 0.91 14.69 0.91 14.69 1 14.35 1 14.35 0.91 12.45 0.91 12.45 1 12.11 1 12.11 0.91 10.155 0.91 10.155 1.525 9.925 1.525  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_4
