# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai32_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai32_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 24.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.67 2.27 13.055 2.27 13.055 2.71 9.67 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.08 2.215 1.31 2.215 1.31 2.785 4.245 2.785 4.245 2.27 7.13 2.27 7.13 2.785 8.78 2.785 8.78 2.215 9.01 2.215 9.01 3.015 6.87 3.015 6.87 2.5 4.475 2.5 4.475 3.015 1.08 3.015  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.37 1.81 7.43 1.81 7.43 1.77 7.69 1.77 7.69 2.555 7.43 2.555 7.43 2.04 3.6 2.04 3.6 2.555 3.37 2.555  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 17.275 1.81 20.31 1.81 20.31 1.77 20.57 1.77 20.57 2.27 20.785 2.27 20.785 2.5 20.31 2.5 20.31 2.04 17.615 2.04 17.615 2.5 17.275 2.5  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 15.035 2.27 15.535 2.27 15.535 2.73 17.845 2.73 17.845 2.27 18.86 2.27 18.86 2.73 22.36 2.73 22.36 2.215 22.59 2.215 22.59 2.96 18.89 2.96 18.89 3.27 18.63 3.27 18.63 2.5 18.075 2.5 18.075 2.96 15.305 2.96 15.305 2.5 15.035 2.5  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.467 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.53 3.09 15.115 3.09 15.115 3.19 16.93 3.19 16.93 3.45 17.21 3.45 17.21 3.77 21.08 3.77 21.08 3.19 22.82 3.19 22.82 1.565 20.675 1.565 20.675 1.54 20.07 1.54 20.07 1.57 15.53 1.57 15.53 1.14 15.76 1.14 15.76 1.34 17.77 1.34 17.77 1.14 18 1.14 18 1.34 19.955 1.34 19.955 1.14 20.78 1.14 20.78 1.335 22.25 1.335 22.25 1.14 23.05 1.14 23.05 3.42 21.31 3.42 21.31 4 16.7 4 16.7 3.42 14.925 3.42 14.925 3.32 12.8 3.32 12.8 3.9 12.57 3.9 12.57 3.32 10.76 3.32 10.76 3.9 10.53 3.9  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 2.59 4.59 2.59 3.705 2.82 3.705 2.82 4.59 7.07 4.59 7.07 3.705 7.3 3.705 7.3 4.59 14.02 4.59 14.51 4.59 14.51 3.56 14.74 3.56 14.74 4.59 18.84 4.59 18.84 4.345 19.07 4.345 19.07 4.59 23.28 4.59 23.28 3.09 23.51 3.09 23.51 4.59 23.6 4.59 24.08 4.59 24.08 5.49 23.6 5.49 14.02 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 24.08 -0.45 24.08 0.45 13 0.45 13 1.11 12.77 1.11 12.77 0.45 10.76 0.45 10.76 1.11 10.53 1.11 10.53 0.45 8.52 0.45 8.52 1.11 8.29 1.11 8.29 0.45 6.28 0.45 6.28 1.11 6.05 1.11 6.05 0.45 4.04 0.45 4.04 1.11 3.81 1.11 3.81 0.45 1.8 0.45 1.8 1.11 1.57 1.11 1.57 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.5 3.09 0.73 3.09 0.73 3.245 4.88 3.245 4.88 3.09 5.11 3.09 5.11 3.245 7.76 3.245 7.76 4.13 11.55 4.13 11.55 3.55 11.78 3.55 11.78 4.13 13.79 4.13 13.79 3.55 14.02 3.55 14.02 4.36 7.53 4.36 7.53 3.475 5.11 3.475 5.11 3.9 4.88 3.9 4.88 3.475 0.73 3.475 0.73 3.9 0.5 3.9  ;
        POLYGON 0.45 0.77 0.68 0.77 0.68 1.35 2.69 1.35 2.69 0.77 2.92 0.77 2.92 1.35 4.93 1.35 4.93 0.77 5.16 0.77 5.16 1.35 7.17 1.35 7.17 0.73 7.4 0.73 7.4 1.31 7.95 1.31 7.95 1.35 9.41 1.35 9.41 0.77 9.64 0.77 9.64 1.35 11.65 1.35 11.65 0.77 11.88 0.77 11.88 1.35 13.89 1.35 13.89 0.68 23.6 0.68 23.6 1.58 23.37 1.58 23.37 0.91 21.36 0.91 21.36 1.105 21.13 1.105 21.13 0.91 19.12 0.91 19.12 1.11 18.89 1.11 18.89 0.91 16.88 0.91 16.88 1.11 16.65 1.11 16.65 0.91 14.12 0.91 14.12 1.58 7.82 1.58 7.82 1.54 7.3 1.54 7.3 1.58 0.45 1.58  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai32_4
