# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.79 1.87 2.55 1.87 2.55 2.5 3.185 2.5 4.07 2.5 4.07 1.77 4.355 1.77 4.355 2.73 3.185 2.73 2.32 2.73 2.32 2.1 1.79 2.1  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.77 2.235 1.46 2.235 1.46 2.33 2.09 2.33 2.09 2.96 3.185 2.96 5.145 2.96 5.145 2.18 5.375 2.18 5.375 3.19 3.185 3.19 1.86 3.19 1.86 2.71 1.27 2.71 1.27 2.465 0.77 2.465  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER METAL1 ;
        POLYGON 7.43 1.21 7.665 1.21 7.665 0.84 7.895 0.84 7.895 4.23 7.665 4.23 7.665 1.59 7.43 1.59  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.585 0.475 3.585 0.475 4.59 2.285 4.59 2.285 3.585 2.515 3.585 2.515 4.59 3.185 4.59 5.725 4.59 5.725 3.88 5.955 3.88 5.955 4.59 6.645 4.59 6.645 3.585 6.875 3.585 6.875 4.59 7.37 4.59 8.685 4.59 8.685 3.585 8.915 3.585 8.915 4.59 9.52 4.59 9.52 5.49 7.37 5.49 3.185 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 9.015 0.45 9.015 1.65 8.785 1.65 8.785 0.45 6.775 0.45 6.775 1.445 6.545 1.445 6.545 0.45 2.515 0.45 2.515 1.18 2.285 1.18 2.285 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.84 0.475 0.84 0.475 1.41 3.185 1.41 3.185 2.27 2.955 2.27 2.955 1.64 0.475 1.64 0.475 2.94 1.495 2.94 1.495 4.31 1.265 4.31 1.265 3.17 0.245 3.17  ;
        POLYGON 3.585 0.68 6.055 0.68 6.055 1.49 5.825 1.49 5.825 0.91 3.815 0.91 3.815 1.65 3.585 1.65  ;
        POLYGON 3.685 3.42 5.605 3.42 5.605 1.95 4.705 1.95 4.705 1.14 4.935 1.14 4.935 1.72 5.825 1.72 5.825 1.88 7.37 1.88 7.37 2.11 5.835 2.11 5.835 3.65 3.915 3.65 3.915 4.23 3.685 4.23  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_2
