# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.06 2.27 3.51 2.27 3.51 1.77 3.77 1.77 3.77 1.81 4.84 1.81 4.84 2.27 6.57 2.27 6.57 2.5 4.61 2.5 4.61 2.04 3.77 2.04 3.77 2.5 3.06 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.25 2.27 2.83 2.27 2.83 2.73 4.04 2.73 4.04 2.27 4.38 2.27 4.38 2.73 6.8 2.73 6.8 2.27 8.81 2.27 8.81 2.5 7.03 2.5 7.03 2.96 2.6 2.96 2.6 2.5 1.25 2.5  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.27 2.27 11.35 2.27 11.35 1.77 11.61 1.77 11.61 2.27 12.85 2.27 12.85 2.5 10.27 2.5  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.7986 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.02 3.19 12.745 3.19 12.745 4.36 12.515 4.36 12.515 3.42 10.555 3.42 10.555 4.36 10.325 4.36 10.325 3.42 7.145 3.42 7.145 4.36 6.915 4.36 6.915 3.42 2.715 3.42 2.715 4.36 2.485 4.36 2.485 3.42 0.79 3.42 0.79 1.81 1.365 1.81 1.365 1.14 1.595 1.14 1.595 1.81 2.95 1.81 2.95 1.14 4.12 1.14 4.12 1.34 5.845 1.34 5.845 1.14 6.075 1.14 6.075 1.34 8.085 1.34 8.085 1.14 8.315 1.14 8.315 1.57 3.935 1.57 3.935 1.48 3.21 1.48 3.21 2.04 1.02 2.04  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.65 0.575 3.65 0.575 4.59 4.675 4.59 4.675 3.65 4.905 3.65 4.905 4.59 9.105 4.59 9.105 3.65 9.335 3.65 9.335 4.59 11.345 4.59 11.345 3.65 11.575 3.65 11.575 4.59 13.635 4.59 13.635 3.65 13.865 3.65 13.865 4.59 13.915 4.59 14.56 4.59 14.56 5.49 13.915 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 12.795 0.45 12.795 1.11 12.565 1.11 12.565 0.45 10.555 0.45 10.555 1.195 10.325 1.195 10.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 9.435 0.68 9.435 1.425 10.95 1.425 10.95 1.31 11.445 1.31 11.445 0.73 11.905 0.73 11.905 1.35 13.685 1.35 13.685 0.77 13.915 0.77 13.915 1.58 11.775 1.58 11.775 1.54 11.15 1.54 11.15 1.655 9.205 1.655 9.205 0.91 7.195 0.91 7.195 1.11 6.965 1.11 6.965 0.91 4.955 0.91 4.955 1.11 4.725 1.11 4.725 0.91 2.715 0.91 2.715 1.58 2.485 1.58 2.485 0.91 0.475 0.91 0.475 1.58 0.245 1.58  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_4
