# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 3.36 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.015 1.77 1.015 2.71 0.71 2.71  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 2.89 2.665 2.89 2.665 1.59 2.39 1.59 2.39 0.74 2.895 0.74 2.895 3.775 2.39 3.775  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.4 1.595 3.4 1.595 4.59 2.215 4.59 3.36 4.59 3.36 5.49 2.215 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 3.36 -0.45 3.36 0.45 1.595 0.45 1.595 1.08 1.365 1.08 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.93 2.94 1.93 1.54 0.245 1.54 0.245 0.74 0.475 0.74 0.475 1.31 2.16 1.31 2.16 1.775 2.215 1.775 2.215 2.585 2.16 2.585 2.16 3.17 0.575 3.17 0.575 3.775 0.345 3.775  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_1
