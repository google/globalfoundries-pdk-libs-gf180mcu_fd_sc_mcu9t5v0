# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.68 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.63 1.21 4.89 1.21 4.89 2.115 4.63 2.115  ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.235 1.575 2.235 1.575 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.71 2.33 14.885 2.33 14.885 0.845 15.115 0.845 15.115 3.685 14.71 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.895 1.595 3.895 1.595 4.59 3.185 4.59 3.185 3.905 3.415 3.905 3.415 4.59 6.115 4.59 7.205 4.59 7.205 3.045 7.435 3.045 7.435 4.59 7.875 4.59 8.855 4.59 12.025 4.59 12.025 3.145 12.255 3.145 12.255 4.59 12.75 4.59 13.765 4.59 13.765 3.875 13.995 3.875 13.995 4.59 14.49 4.59 15.68 4.59 15.68 5.49 14.49 5.49 12.75 5.49 8.855 5.49 7.875 5.49 6.115 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 15.68 -0.45 15.68 0.45 13.995 0.45 13.995 1.165 13.765 1.165 13.765 0.45 12.155 0.45 12.155 1.265 11.925 1.265 11.925 0.45 7.525 0.45 7.525 0.625 7.295 0.625 7.295 0.45 3.435 0.45 3.435 1.435 3.205 1.435 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 3.425 1.805 3.425 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.445 6.115 3.445 6.115 4.315 5.885 4.315 5.885 3.675 1.94 3.675 1.94 3.655 0.575 3.655 0.575 4.235 0.345 4.235  ;
        POLYGON 5.165 1.315 5.395 1.315 5.395 2.415 7.875 2.415 7.875 2.755 5.395 2.755 5.395 3.215 5.165 3.215  ;
        POLYGON 6.685 1.775 8.225 1.775 8.225 1.315 8.855 1.315 8.855 1.655 8.455 1.655 8.455 3.685 8.225 3.685 8.225 2.115 6.685 2.115  ;
        POLYGON 2.385 2.525 3.845 2.525 3.845 1.895 2.485 1.895 2.485 1.315 2.715 1.315 2.715 1.665 3.845 1.665 3.845 0.69 5.89 0.69 5.89 0.855 9.01 0.855 9.01 0.69 10.735 0.69 10.735 2.755 10.505 2.755 10.505 1.085 5.665 1.085 5.665 0.92 4.075 0.92 4.075 2.755 2.615 2.755 2.615 3.215 2.385 3.215  ;
        POLYGON 9.745 1.315 9.975 1.315 9.975 3.455 11.565 3.455 11.565 2.47 12.75 2.47 12.75 2.7 11.795 2.7 11.795 3.685 9.745 3.685  ;
        POLYGON 11.265 1.775 13.045 1.775 13.045 1.315 13.275 1.315 13.275 1.83 14.49 1.83 14.49 2.06 13.275 2.06 13.275 3.685 13.045 3.685 13.045 2.115 11.265 2.115  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffq_1
