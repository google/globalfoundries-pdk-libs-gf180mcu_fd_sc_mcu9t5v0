# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 23.52 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.945 2.33 4.03 2.33 4.03 2.71 2.945 2.71  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER METAL1 ;
        POLYGON 13.53 2.22 14.515 2.22 14.515 2.71 13.53 2.71  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.24 1.57 2.24 1.57 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER METAL1 ;
        POLYGON 19.11 2.875 20.92 2.875 21.59 2.875 21.59 1.655 19.405 1.655 19.405 0.845 19.64 0.845 19.64 1.395 21.59 1.395 21.59 0.845 21.88 0.845 21.88 3.685 21.15 3.685 21.15 3.105 20.92 3.105 19.34 3.105 19.34 3.685 19.11 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.09 4.59 3.305 4.59 3.305 3.615 3.535 3.615 3.535 4.59 5.295 4.59 7.51 4.59 7.51 3.615 7.74 3.615 7.74 4.59 9.715 4.59 9.715 3.885 10.055 3.885 10.055 4.59 11.38 4.59 13.79 4.59 13.79 3.515 14.02 3.515 14.02 4.59 15.04 4.59 15.83 4.59 15.83 3.045 16.06 3.045 16.06 4.59 18.09 4.59 18.09 3.875 18.32 3.875 18.32 4.59 20.13 4.59 20.13 3.875 20.36 3.875 20.36 4.59 20.92 4.59 22.17 4.59 22.17 3.875 22.4 3.875 22.4 4.59 23.52 4.59 23.52 5.49 20.92 5.49 15.04 5.49 11.38 5.49 5.295 5.49 2.09 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 23.52 -0.45 23.52 0.45 23 0.45 23 1.165 22.77 1.165 22.77 0.45 20.76 0.45 20.76 1.165 20.53 1.165 20.53 0.45 18.52 0.45 18.52 1.165 18.29 1.165 18.29 0.45 16.335 0.45 16.335 0.64 15.995 0.64 15.995 0.45 7.795 0.45 7.795 1.37 7.455 1.37 7.455 0.45 3.435 0.45 3.435 1.425 3.205 1.425 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 2.94 1.86 2.94 1.86 1.685 0.245 1.685 0.245 1.315 0.475 1.315 0.475 1.455 2.09 1.455 2.09 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.325 1.315 4.555 1.315 4.555 3.785 4.325 3.785  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 3.155 3.995 3.155 3.995 4.13 5.295 4.13 5.295 4.36 3.765 4.36 3.765 3.385 2.615 3.385 2.615 3.685 2.385 3.685  ;
        POLYGON 5.445 1.315 5.675 1.315 5.675 2.29 6.565 2.29 6.565 2.11 8.235 2.11 8.235 2.34 6.79 2.34 6.79 2.52 5.82 2.52 5.82 3.785 5.445 3.785  ;
        POLYGON 6 1.65 9.09 1.65 9.09 0.68 10.315 0.68 10.315 0.91 9.32 0.91 9.32 1.88 6.34 1.88 6.34 2.06 6 2.06  ;
        POLYGON 7.015 2.57 9.55 2.57 9.55 1.315 9.78 1.315 9.78 2.57 10.995 2.57 10.995 3.16 10.655 3.16 10.655 2.8 8.815 2.8 8.815 3.26 8.475 3.26 8.475 2.8 7.015 2.8  ;
        POLYGON 6.115 3.155 8.2 3.155 8.2 3.49 9.32 3.49 9.32 3.425 11.38 3.425 11.38 4.315 11.15 4.315 11.15 3.655 9.545 3.655 9.545 3.72 7.97 3.72 7.97 3.385 6.455 3.385 6.455 4.36 6.115 4.36  ;
        POLYGON 13.3 2.985 14.81 2.985 14.81 2.875 15.04 2.875 15.04 3.685 14.81 3.685 14.81 3.215 13.07 3.215 13.07 1.655 11.83 1.655 11.83 1.315 14.1 1.315 14.1 1.655 13.3 1.655  ;
        POLYGON 10.71 0.855 15.91 0.855 15.91 1.83 16.775 1.83 16.775 2.06 15.68 2.06 15.68 1.085 11.6 1.085 11.6 1.885 11.96 1.885 11.96 3.685 11.73 3.685 11.73 2.115 11.37 2.115 11.37 1.425 10.71 1.425  ;
        POLYGON 15.25 2.18 15.48 2.18 15.48 2.29 17.075 2.29 17.075 0.845 17.4 0.845 17.4 2.03 20.92 2.03 20.92 2.325 17.305 2.325 17.305 3.685 17.07 3.685 17.07 2.52 15.25 2.52  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffsnq_4
