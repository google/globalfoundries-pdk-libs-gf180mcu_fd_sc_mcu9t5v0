* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
*.PININFO I0:I I1:I I2:I I3:I S0:I S1:I Z:O VDD:P VNW:P VPW:P VSS:G
*.EQN Z=((S0 * ((S1 * I3) + (!S1 * I1))) + (!S0 * ((S1 * I2) + (!S1 * I0))))
M_MN5 int01 I2 VSS VPW nfet_05v0 W=0.660000U L=0.600000U
M_MN9 int02 sel1_n int01 VPW nfet_05v0 W=0.660000U L=0.600000U
M_MN10 int07 S0 int02 VPW nfet_05v0 W=0.660000U L=0.600000U
M_MN6 VSS I3 int07 VPW nfet_05v0 W=0.660000U L=0.600000U
M_instance_22 Z int03 VSS VPW nfet_05v0 W=0.900000U L=0.600000U
M_MN12 int03 S1 int02 VPW nfet_05v0 W=0.660000U L=0.600000U
M_MN11 int04 sel2_n int03 VPW nfet_05v0 W=0.660000U L=0.600000U
M_MN2 VSS S1 sel2_n VPW nfet_05v0 W=0.660000U L=0.600000U
M_MN4 int06 I1 VSS VPW nfet_05v0 W=0.660000U L=0.600000U
M_MN8 int04 S0 int06 VPW nfet_05v0 W=0.660000U L=0.600000U
M_MN7 int05 sel1_n int04 VPW nfet_05v0 W=0.660000U L=0.600000U
M_MN3 VSS I0 int05 VPW nfet_05v0 W=0.660000U L=0.600000U
M_MN1 sel1_n S0 VSS VPW nfet_05v0 W=0.660000U L=0.600000U
M_MP2 int01 I2 VDD VNW pfet_05v0 W=0.915000U L=0.500000U
M_MP9 int02 S0 int01 VNW pfet_05v0 W=0.915000U L=0.500000U
M_MP10 int07 sel1_n int02 VNW pfet_05v0 W=0.915000U L=0.500000U
M_MP6 VDD I3 int07 VNW pfet_05v0 W=0.915000U L=0.500000U
M_instance_1 Z int03 VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_MP12 int03 sel2_n int02 VNW pfet_05v0 W=0.915000U L=0.500000U
M_MP11 int04 S1 int03 VNW pfet_05v0 W=0.915000U L=0.500000U
M_MP5 VDD S1 sel2_n VNW pfet_05v0 W=0.915000U L=0.500000U
M_MP4 int06 I1 VDD VNW pfet_05v0 W=0.915000U L=0.500000U
M_MP8 int04 sel1_n int06 VNW pfet_05v0 W=0.915000U L=0.500000U
M_MP7 int05 S0 int04 VNW pfet_05v0 W=0.915000U L=0.500000U
M_MP3 VDD I0 int05 VNW pfet_05v0 W=0.915000U L=0.500000U
M_MP1 sel1_n S0 VDD VNW pfet_05v0 W=0.915000U L=0.500000U
.ENDS
