# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.19 1.21 19.45 1.21 19.45 2.03 19.19 2.03  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.83 2.15 16.09 2.15 16.09 2.71 15.83 2.71  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.7 2.33 1.08 2.33 1.08 2.71 0.7 2.71  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.12 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 2.15 4.89 2.15 4.89 2.71 4.63 2.71  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.36 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.35 1.77 3.885 1.77 3.885 2.22 2.58 2.22 2.58 2.71 2.35 2.71  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.24 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.79 1.945 12.47 1.945 12.47 1.21 12.73 1.21 12.73 1.945 13.135 1.945 13.135 2.83 12.905 2.83 12.905 2.175 11.79 2.175  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1632 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.59 1.23 6.82 1.23 6.82 1.8 8.83 1.8 8.83 1.21 9.37 1.21 9.37 3.38 9.075 3.38 9.075 2.03 6.825 2.03 6.825 3.38 6.59 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.41 4.59 0.41 3.04 0.64 3.04 0.64 4.59 1.66 4.59 5.355 4.59 5.355 4.07 5.585 4.07 5.585 4.59 7.835 4.59 7.835 4.07 8.065 4.07 8.065 4.59 10.095 4.59 10.095 3.44 10.325 3.44 10.325 4.59 11.655 4.59 12.675 4.59 15.245 4.59 15.245 3.4 15.475 3.4 15.475 4.59 17.675 4.59 19.585 4.59 19.585 3.04 19.815 3.04 19.815 4.59 21.035 4.59 21.28 4.59 21.28 5.49 21.035 5.49 17.675 5.49 12.675 5.49 11.655 5.49 1.66 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 19.915 0.45 19.915 1.57 19.685 1.57 19.685 0.45 15.435 0.45 15.435 1.57 15.205 1.57 15.205 0.45 10.18 0.45 10.18 1.57 9.95 1.57 9.95 0.45 7.94 0.45 7.94 1.57 7.71 1.57 7.71 0.45 5.7 0.45 5.7 1.57 5.47 1.57 5.47 0.45 0.54 0.45 0.54 1.57 0.31 1.57 0.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.43 1.23 1.66 1.23 1.66 3.85 1.43 3.85  ;
        POLYGON 4.115 1.695 4.35 1.695 4.35 1.23 4.58 1.23 4.58 1.925 4.345 1.925 4.345 3.38 4.115 3.38  ;
        POLYGON 2.12 3.61 2.79 3.61 2.79 3.04 3.02 3.04 3.02 3.61 9.635 3.61 9.635 2.98 10.87 2.98 10.87 1.23 11.1 1.23 11.1 3.04 11.655 3.04 11.655 3.85 11.425 3.85 11.425 3.27 10.945 3.27 10.945 3.21 9.865 3.21 9.865 3.84 3.02 3.84 3.02 3.85 1.89 3.85 1.89 1.285 3.515 1.285 3.515 1.515 2.12 1.515  ;
        POLYGON 11.56 2.405 12.675 2.405 12.675 3.85 12.445 3.85 12.445 2.635 11.33 2.635 11.33 1 10.64 1 10.64 2.03 9.885 2.03 9.885 2.71 9.655 2.71 9.655 1.8 10.41 1.8 10.41 0.77 12.235 0.77 12.235 1.57 12.005 1.57 12.005 1 11.56 1  ;
        POLYGON 13.925 1.23 14.455 1.23 14.455 3.85 13.925 3.85  ;
        POLYGON 16.325 1.23 16.555 1.23 16.555 3.85 16.325 3.85  ;
        POLYGON 13.125 1.23 13.695 1.23 13.695 4.08 14.785 4.08 14.785 2.94 15.935 2.94 15.935 4.08 17.445 4.08 17.445 1.23 17.675 1.23 17.675 4.31 15.705 4.31 15.705 3.17 15.015 3.17 15.015 4.31 13.465 4.31 13.465 1.57 13.125 1.57  ;
        POLYGON 17.945 1.285 18.85 1.285 18.85 1.515 18.175 1.515 18.175 2.72 18.795 2.72 18.795 3.85 18.565 3.85 18.565 2.95 17.945 2.95  ;
        POLYGON 18.405 2.15 18.635 2.15 18.635 2.26 20.805 2.26 20.805 1.23 21.035 1.23 21.035 3.85 20.705 3.85 20.705 2.49 18.405 2.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_4
