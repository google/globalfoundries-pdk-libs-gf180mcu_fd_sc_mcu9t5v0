# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.64 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 7.99 1.21 8.25 1.21 8.25 1.83 8.645 1.83 8.645 2.15 7.99 2.15  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.13 1.77 6.01 1.77 6.01 2.15 5.13 2.15  ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.3 1.775 6.53 1.775 6.53 2.47 9.05 2.47 9.05 1.83 9.665 1.83 9.665 2.06 9.43 2.06 9.43 2.7 6.3 2.7  ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.5505 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.42 0.68 1.65 0.68 1.65 2.33 3.66 2.33 3.66 0.68 3.89 0.68 3.89 4.36 3.61 4.36 3.61 2.71 1.65 2.71 1.65 4.36 1.42 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.35 4.59 0.35 3.55 0.58 3.55 0.58 4.59 2.49 4.59 2.49 3.55 2.72 3.55 2.72 4.59 4.68 4.59 4.68 3.55 4.91 3.55 4.91 4.59 7.41 4.59 8.94 4.59 8.94 3.55 9.17 3.55 9.17 4.59 10.29 4.59 10.64 4.59 10.64 5.49 10.29 5.49 7.41 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 10.64 -0.45 10.64 0.45 9.17 0.45 9.17 1.02 8.94 1.02 8.94 0.45 5.01 0.45 5.01 1.02 4.78 1.02 4.78 0.45 2.77 0.45 2.77 1.49 2.54 1.49 2.54 0.45 0.53 0.45 0.53 1.49 0.3 1.49 0.3 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 4.9 2.93 7.41 2.93 7.41 4.36 7.18 4.36 7.18 3.16 4.67 3.16 4.67 2.115 4.24 2.115 4.24 1.775 4.67 1.775 4.67 1.31 6.74 1.31 6.74 0.68 6.97 0.68 6.97 1.54 4.9 1.54  ;
        POLYGON 7.125 1.83 7.53 1.83 7.53 0.75 8.71 0.75 8.71 1.25 10.06 1.25 10.06 0.68 10.29 0.68 10.29 4.36 9.96 4.36 9.96 1.48 8.48 1.48 8.48 0.98 7.76 0.98 7.76 2.06 7.125 2.06  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_4
