* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__xnor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(!((!((A1 * A2) + !(A1 + A2)) * A3) + !(!((A1 * A2) + !(A1 + A2)) + A3)))
M_i_14 I A2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_15 VSS A1 I VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 I2 I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_0 net_0 A1 I2 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_18 I3 I2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_19 VSS A3 I3 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_10 Z_neg I3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8 net_2 A3 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9 VSS I2 net_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_3 VSS Z_neg ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_2 ZN Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_1 VSS Z_neg ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_0 ZN Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_16 net_4 A2 I VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_17 VDD A1 net_4 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_5 net_1 I VDD VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_3 I2 A1 net_1 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_4 net_1 A2 I2 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_20 net_5 I2 I3 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_21 VDD A3 net_5 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_13 net_3 I3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11 Z_neg A3 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_12 net_3 I2 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 VDD Z_neg ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 ZN Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 VDD Z_neg ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 ZN Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
