# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.868 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.06 2.27 3.58 2.27 3.58 1.77 4.89 1.77 4.89 2.27 6.62 2.27 6.62 2.5 4.63 2.5 4.63 2 3.81 2 3.81 2.5 3.06 2.5  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.868 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.2 2.27 2.83 2.27 2.83 2.73 4.04 2.73 4.04 2.27 4.38 2.27 4.38 2.73 6.85 2.73 6.85 2.27 8.86 2.27 8.86 2.5 7.08 2.5 7.08 2.96 2.6 2.96 2.6 2.5 1.2 2.5  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.0913 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.26 1.365 1.26 1.365 0.68 1.595 0.68 1.595 1.26 3.605 1.26 3.605 0.68 3.835 0.68 3.835 1.26 5.845 1.26 5.845 0.68 6.075 0.68 6.075 1.26 8.085 1.26 8.085 0.68 8.315 0.68 8.315 1.49 0.97 1.49 0.97 3.19 7.145 3.19 7.145 4.36 6.915 4.36 6.915 3.42 2.715 3.42 2.715 4.36 2.485 4.36 2.485 3.42 0.71 3.42  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.65 0.525 3.65 0.525 4.59 4.675 4.59 4.675 3.65 4.905 3.65 4.905 4.59 9.155 4.59 9.155 3.65 9.385 3.65 9.385 4.59 10.08 4.59 10.08 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 9.435 0.45 9.435 1.4 9.205 1.4 9.205 0.45 7.195 0.45 7.195 1.02 6.965 1.02 6.965 0.45 4.955 0.45 4.955 1.02 4.725 1.02 4.725 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor2_4
