# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 22.4 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.77 4.33 1.77 4.33 2.225 4.835 2.225 4.835 2.71 4.07 2.71  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.41 1.77 0.41 2.225 1.015 2.225 1.015 2.71 0.15 2.71  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.77 2.135 1.77 2.135 2.71 1.83 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 1.77 7.69 1.77 7.69 2.71 7.43 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.70205 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.79 0.845 21.13 0.845 21.13 4.25 20.79 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.44 1.595 3.44 1.595 4.59 2.895 4.59 5.235 4.59 5.235 3.905 5.465 3.905 5.465 4.59 7.83 4.59 7.83 3.905 8.17 3.905 8.17 4.59 10.685 4.59 11.125 4.59 13.235 4.59 13.235 3.44 13.465 3.44 13.465 4.59 14.485 4.59 17.645 4.59 17.645 3.6 17.875 3.6 17.875 4.59 18.37 4.59 19.41 4.59 19.735 4.59 19.735 3.88 19.965 3.88 19.965 4.59 21.81 4.59 21.81 3.88 22.04 3.88 22.04 4.59 22.4 4.59 22.4 5.49 19.41 5.49 18.37 5.49 14.485 5.49 11.125 5.49 10.685 5.49 2.895 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 22.4 -0.45 22.4 0.45 22.155 0.45 22.155 1.165 21.925 1.165 21.925 0.45 19.915 0.45 19.915 1.6 19.685 1.6 19.685 0.45 17.975 0.45 17.975 1.59 17.745 1.59 17.745 0.45 13.1 0.45 13.1 0.62 12.87 0.62 12.87 0.45 7.795 0.45 7.795 0.62 7.565 0.62 7.565 0.45 5.735 0.45 5.735 0.62 5.505 0.62 5.505 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.98 2.665 2.98 2.665 1.54 0.245 1.54 0.245 0.79 0.475 0.79 0.475 1.31 2.895 1.31 2.895 3.21 0.575 3.21 0.575 4.25 0.345 4.25  ;
        POLYGON 6.865 2.875 7.095 2.875 7.095 2.985 8.325 2.985 8.325 1.54 6.455 1.54 6.455 1.65 6.225 1.65 6.225 1.31 8.555 1.31 8.555 3.215 6.865 3.215  ;
        POLYGON 3.325 0.79 3.555 0.79 3.555 0.85 9.855 0.85 9.855 1.43 9.625 1.43 9.625 1.08 3.555 1.08 3.555 1.13 3.325 1.13  ;
        POLYGON 3.375 3.44 3.605 3.44 3.605 4.02 4.775 4.02 4.775 3.445 10.685 3.445 10.685 3.785 10.455 3.785 10.455 3.675 5.005 3.675 5.005 4.25 3.375 4.25  ;
        POLYGON 8.905 1.31 9.135 1.31 9.135 2.225 11.125 2.225 11.125 2.565 9.135 2.565 9.135 3.215 8.905 3.215  ;
        POLYGON 10.745 1.31 11.705 1.31 11.705 1.765 13.755 1.765 13.755 2.565 13.525 2.565 13.525 1.995 11.705 1.995 11.705 4.25 11.475 4.25 11.475 1.65 10.745 1.65  ;
        POLYGON 12.795 2.225 13.025 2.225 13.025 2.795 14.205 2.795 14.205 1.31 14.485 1.31 14.485 4.25 14.255 4.25 14.255 3.025 12.795 3.025  ;
        POLYGON 11.37 0.685 11.71 0.685 11.71 0.85 14.73 0.85 14.73 0.685 16.015 0.685 16.015 2.91 15.785 2.91 15.785 1.08 11.37 1.08  ;
        POLYGON 15.325 1.31 15.555 1.31 15.555 3.14 17.665 3.14 17.665 2.28 18.37 2.28 18.37 2.51 17.895 2.51 17.895 3.37 15.555 3.37 15.555 4.25 15.325 4.25  ;
        POLYGON 17.205 1.82 18.865 1.82 18.865 0.79 19.095 0.79 19.095 2.225 19.41 2.225 19.41 2.565 18.895 2.565 18.895 4.25 18.665 4.25 18.665 2.05 17.435 2.05 17.435 2.565 17.205 2.565  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_2
