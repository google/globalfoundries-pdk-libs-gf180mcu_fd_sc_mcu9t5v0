# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 1.21 4.89 1.21 4.89 2.52 4.63 2.52  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.41 1.77 0.41 2.18 0.915 2.18 0.915 2.71 0.15 2.71  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.848 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 1.77 1.53 1.77 1.53 2.18 2.02 2.18 2.02 2.71 1.27 2.71  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 1.77 6.835 1.77 6.835 2.71 6.31 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.19 1.21 19.445 1.21 19.445 0.79 19.725 0.79 19.725 3.69 19.495 3.69 19.495 2.71 19.19 2.71  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.315 4.59 1.315 3.44 1.545 3.44 1.545 4.59 2.775 4.59 5.03 4.59 5.03 3.965 5.37 3.965 5.37 4.59 7.18 4.59 7.18 3.995 7.52 3.995 7.52 4.59 9.845 4.59 10.285 4.59 12.595 4.59 12.595 3.44 12.825 3.44 12.825 4.59 14.375 4.59 17.025 4.59 17.025 3.595 17.255 3.595 17.255 4.59 17.93 4.59 18.955 4.59 20.515 4.59 20.515 3.88 20.745 3.88 20.745 4.59 21.28 4.59 21.28 5.49 18.955 5.49 17.93 5.49 14.375 5.49 10.285 5.49 9.845 5.49 2.775 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.795 0.45 20.795 1.6 20.565 1.6 20.565 0.45 17.615 0.45 17.615 0.72 17.385 0.72 17.385 0.45 13.15 0.45 13.15 0.505 12.81 0.505 12.81 0.45 7.79 0.45 7.79 0.51 7.45 0.51 7.45 0.45 5.79 0.45 5.79 0.51 5.45 0.51 5.45 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.295 2.98 2.545 2.98 2.545 1.535 0.245 1.535 0.245 0.79 0.475 0.79 0.475 1.305 2.775 1.305 2.775 3.21 0.525 3.21 0.525 4.25 0.295 4.25  ;
        POLYGON 6.03 2.935 6.26 2.935 6.26 3.045 8.125 3.045 8.125 1.54 6.165 1.54 6.165 1.2 8.355 1.2 8.355 3.275 6.03 3.275  ;
        POLYGON 3.325 0.74 9.795 0.74 9.795 1.48 9.565 1.48 9.565 0.97 3.555 0.97 3.555 1.13 3.325 1.13  ;
        POLYGON 3.125 3.44 3.355 3.44 3.355 3.505 9.845 3.505 9.845 3.845 9.615 3.845 9.615 3.735 3.355 3.735 3.355 4.25 3.125 4.25  ;
        POLYGON 8.705 1.22 9.075 1.22 9.075 2.18 10.285 2.18 10.285 2.52 8.935 2.52 8.935 3.26 8.705 3.26  ;
        POLYGON 10.685 1.36 10.915 1.36 10.915 1.72 13.665 1.72 13.665 2.52 13.435 2.52 13.435 1.95 10.915 1.95 10.915 4.25 10.685 4.25  ;
        POLYGON 12.205 2.18 12.435 2.18 12.435 2.75 14.145 2.75 14.145 1.36 14.375 1.36 14.375 4.25 14.015 4.25 14.015 2.98 12.205 2.98  ;
        POLYGON 11.365 0.68 11.595 0.68 11.595 0.735 16.065 0.735 16.065 2.905 15.725 2.905 15.725 1.02 11.365 1.02  ;
        POLYGON 15.265 1.36 15.495 1.36 15.495 3.135 17.59 3.135 17.59 2.235 17.93 2.235 17.93 3.365 15.495 3.365 15.495 4.25 15.265 4.25  ;
        POLYGON 18.225 2.29 18.725 2.29 18.725 1.545 16.97 1.545 16.97 2.465 16.63 2.465 16.63 1.315 18.955 1.315 18.955 2.52 18.455 2.52 18.455 4.25 18.225 4.25  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffq_1
