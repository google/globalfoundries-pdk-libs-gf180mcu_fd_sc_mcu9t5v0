# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.795 2.215 2.09 2.215 2.09 2.71 1.795 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 2.27 1.54 2.27 1.54 2.94 2.39 2.94 2.39 2.27 4.33 2.27 4.33 2.71 2.62 2.71 2.62 3.17 1.2 3.17  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.33 2.27 5.67 2.27 5.67 2.94 6.87 2.94 6.87 2.215 8.535 2.215 8.535 3.17 5.33 3.17  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.23 2.27 6.57 2.27 6.57 2.71 6.23 2.71  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.0258 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.97 3.375 1.095 3.375 1.095 4.07 2.435 4.07 2.435 3.4 8.095 3.4 8.095 4.36 7.865 4.36 7.865 3.63 6.055 3.63 6.055 4.36 5.825 4.36 5.825 3.63 2.665 3.63 2.665 4.36 0.865 4.36 0.865 3.58 0.74 3.58 0.74 1.14 1.595 1.14 1.595 1.34 3.89 1.34 3.89 1.57 0.97 1.57  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.86 0.575 3.86 0.575 4.59 4.625 4.59 4.625 3.86 4.855 3.86 4.855 4.59 6.845 4.59 6.845 3.86 7.075 3.86 7.075 4.59 8.885 4.59 8.885 3.86 9.115 3.86 9.115 4.59 9.52 4.59 9.52 5.49 9.115 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 7.075 0.45 7.075 1.525 6.845 1.525 6.845 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 4.955 0.68 4.955 1.755 8.885 1.755 8.885 0.77 9.115 0.77 9.115 1.985 4.725 1.985 4.725 1.11 2.485 1.11 2.485 0.91 0.475 0.91 0.475 1.58 0.245 1.58  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_2
