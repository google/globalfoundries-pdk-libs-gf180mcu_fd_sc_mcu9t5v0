# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__or2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.8 2.27 2.14 2.27 2.14 2.71 1.8 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.87 2.27 1.21 2.27 1.21 2.94 2.39 2.94 2.39 2.215 4.275 2.215 4.275 3.17 0.87 3.17  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.5505 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.085 3.09 7.39 3.09 7.62 3.09 7.62 1.59 5.985 1.59 5.985 0.68 6.215 0.68 6.215 1.21 8.225 1.21 8.225 0.68 8.455 0.68 8.455 1.49 7.85 1.49 7.85 3.09 8.405 3.09 8.405 4.36 8.175 4.36 8.175 3.32 7.39 3.32 6.315 3.32 6.315 4.36 6.085 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 4.965 4.59 4.965 3.55 5.195 3.55 5.195 4.59 7.105 4.59 7.105 3.55 7.335 3.55 7.335 4.59 7.39 4.59 9.245 4.59 9.245 3.55 9.475 3.55 9.475 4.59 10.08 4.59 10.08 5.49 7.39 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 9.575 0.45 9.575 1.49 9.345 1.49 9.345 0.45 7.335 0.45 7.335 0.98 7.105 0.98 7.105 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 2.535 3.4 4.505 3.4 4.505 1.97 1.365 1.97 1.365 0.68 1.595 0.68 1.595 1.74 3.605 1.74 3.605 0.68 3.835 0.68 3.835 1.74 4.735 1.74 4.735 2.27 7.39 2.27 7.39 2.5 4.735 2.5 4.735 3.63 2.765 3.63 2.765 4.36 2.535 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or2_4
