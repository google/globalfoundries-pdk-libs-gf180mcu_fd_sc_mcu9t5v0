# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__or3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__or3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.32 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.09 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.92 2.27 3.26 2.27 3.26 2.71 2.92 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.09 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.77 3.72 1.77 3.72 2.27 5.5 2.27 5.5 2.5 3.49 2.5 3.49 2 2.17 2 2.17 2.5 1.83 2.5  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.09 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.27 1.07 2.27 1.07 2.94 6.23 2.94 6.23 2.27 6.57 2.27 6.57 3.17 0.71 3.17  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.459 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.315 3.4 9.67 3.4 9.9 3.4 9.9 1.59 8.265 1.59 8.265 0.68 8.495 0.68 8.495 1.21 10.505 1.21 10.505 0.68 10.735 0.68 10.735 1.49 10.13 1.49 10.13 3.4 10.685 3.4 10.685 4.36 10.455 4.36 10.455 3.63 9.67 3.63 8.545 3.63 8.545 4.36 8.315 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.86 0.575 3.86 0.575 4.59 6.865 4.59 6.865 3.86 7.095 3.86 7.095 4.59 9.335 4.59 9.335 3.86 9.565 3.86 9.565 4.59 9.67 4.59 11.525 4.59 11.525 3.86 11.755 3.86 11.755 4.59 12.32 4.59 12.32 5.49 9.67 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 12.32 -0.45 12.32 0.45 11.855 0.45 11.855 1.385 11.625 1.385 11.625 0.45 9.615 0.45 9.615 0.915 9.385 0.915 9.385 0.45 7.195 0.45 7.195 0.915 6.965 0.915 6.965 0.45 4.955 0.45 4.955 0.915 4.725 0.915 4.725 0.45 2.715 0.45 2.715 0.915 2.485 0.915 2.485 0.45 0.475 0.45 0.475 1.385 0.245 1.385 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 3.655 3.4 6.8 3.4 6.8 1.375 1.365 1.375 1.365 0.68 1.595 0.68 1.595 1.145 3.605 1.145 3.605 0.68 3.835 0.68 3.835 1.145 5.845 1.145 5.845 0.68 6.075 0.68 6.075 1.145 7.03 1.145 7.03 2.27 9.67 2.27 9.67 2.5 7.03 2.5 7.03 3.63 3.885 3.63 3.885 4.36 3.655 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__or3_4
