# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 26.32 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.51 2.33 4.49 2.33 4.49 2.735 3.51 2.735  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.144 ;
    PORT
      LAYER METAL1 ;
        POLYGON 18.63 1.77 18.89 1.77 18.89 2.79 18.63 2.79  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.77 1.175 1.77 1.175 2.735 0.71 2.735  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.77 2.53 1.77 2.53 2.735 1.83 2.735  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.87 1.77 7.4 1.77 7.4 2.735 6.87 2.735  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER METAL1 ;
        POLYGON 22.425 0.84 22.655 0.84 22.655 1.39 24.23 1.39 24.23 1.21 24.665 1.21 24.665 0.84 24.895 0.84 24.895 4.25 24.23 4.25 24.23 1.62 22.655 1.62 22.655 4.25 22.425 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.51 4.59 1.51 3.44 1.74 3.44 1.74 4.59 5.525 4.59 5.525 3.44 5.755 3.44 5.755 4.59 7.64 4.59 7.64 3.94 7.98 3.94 7.98 4.59 9.995 4.59 10.49 4.59 12.825 4.59 12.825 3.45 13.055 3.45 13.055 4.59 14.075 4.59 14.585 4.59 14.585 3.44 14.77 3.44 14.815 3.44 14.815 4.59 15.835 4.59 18.885 4.59 18.885 4.35 19.115 4.35 19.115 4.59 20.595 4.59 20.925 4.59 20.925 3.44 21.085 3.44 21.155 3.44 21.155 4.59 23.495 4.59 23.495 3.44 23.725 3.44 23.725 4.59 25.645 4.59 25.645 3.44 25.875 3.44 25.875 4.59 26.32 4.59 26.32 5.49 21.085 5.49 20.595 5.49 15.835 5.49 14.77 5.49 14.075 5.49 10.49 5.49 9.995 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 26.32 -0.45 26.32 0.45 26.015 0.45 26.015 1.16 25.785 1.16 25.785 0.45 23.775 0.45 23.775 1.16 23.545 1.16 23.545 0.45 21.535 0.45 21.535 1.16 21.305 1.16 21.305 0.45 18.675 0.45 18.675 1.38 18.445 1.38 18.445 0.45 14.175 0.45 14.175 1.38 13.945 1.38 13.945 0.45 8.195 0.45 8.195 0.62 7.965 0.62 7.965 0.45 6.175 0.45 6.175 0.645 5.945 0.645 5.945 0.45 1.815 0.45 1.815 1.08 1.585 1.08 1.585 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.49 2.965 2.985 2.965 2.985 1.54 0.245 1.54 0.245 1.005 0.475 1.005 0.475 1.31 3.215 1.31 3.215 1.87 5.375 1.87 5.375 2.75 5.145 2.75 5.145 2.1 3.215 2.1 3.215 3.195 0.72 3.195 0.72 4.25 0.49 4.25  ;
        POLYGON 6.62 2.965 7.63 2.965 7.63 2.505 8.19 2.505 8.19 1.54 6.57 1.54 6.57 1.31 8.42 1.31 8.42 2.735 7.86 2.735 7.86 3.195 6.62 3.195  ;
        POLYGON 3.765 2.98 6.215 2.98 6.215 3.48 9.765 3.48 9.765 3.44 9.995 3.44 9.995 4.25 9.765 4.25 9.765 3.71 5.985 3.71 5.985 3.21 3.995 3.21 3.995 4.25 3.765 4.25  ;
        POLYGON 3.765 0.875 6.36 0.875 6.36 0.85 8.855 0.85 8.855 0.735 10.255 0.735 10.255 1.38 10.025 1.38 10.025 0.965 9.08 0.965 9.08 1.08 6.465 1.08 6.465 1.105 3.995 1.105 3.995 1.345 3.765 1.345  ;
        POLYGON 8.715 2.505 9.305 2.505 9.305 1.195 9.535 1.195 9.535 2.505 10.49 2.505 10.49 2.735 8.945 2.735 8.945 3.25 8.715 3.25  ;
        POLYGON 11.805 2.99 14.075 2.99 14.075 4.25 13.845 4.25 13.845 3.22 12.035 3.22 12.035 4.25 11.805 4.25  ;
        POLYGON 10.785 2.71 11.145 2.71 11.145 1.07 11.375 1.07 11.375 2.53 14.77 2.53 14.77 2.76 11.37 2.76 11.37 2.94 11.015 2.94 11.015 4.25 10.785 4.25  ;
        POLYGON 12.37 2.07 15.065 2.07 15.065 1.27 15.295 1.27 15.295 3.02 15.835 3.02 15.835 4.25 15.605 4.25 15.605 3.25 15.065 3.25 15.065 2.3 12.37 2.3  ;
        POLYGON 11.67 1.61 14.605 1.61 14.605 0.81 17.095 0.81 17.095 1.84 17.295 1.84 17.295 2.79 17.065 2.79 17.065 2.07 16.865 2.07 16.865 1.04 15.835 1.04 15.835 2.79 15.605 2.79 15.605 1.04 14.835 1.04 14.835 1.84 12.01 1.84 12.01 2.015 11.67 2.015  ;
        POLYGON 17.325 1.27 17.755 1.27 17.755 3.44 17.875 3.44 17.875 3.78 17.525 3.78 17.525 1.61 17.325 1.61  ;
        POLYGON 16.185 1.27 16.415 1.27 16.415 2.885 16.855 2.885 16.855 4.02 18.4 4.02 18.4 3.89 19.375 3.89 19.375 3.93 20.365 3.93 20.365 2.855 20.345 2.855 20.345 2.515 20.595 2.515 20.595 4.16 19.245 4.16 19.245 4.12 18.68 4.12 18.68 4.245 18.45 4.245 18.45 4.25 16.625 4.25 16.625 3.115 16.185 3.115  ;
        POLYGON 18.005 2.45 18.235 2.45 18.235 3.02 19.885 3.02 19.885 1.985 20.585 1.985 20.585 0.8 20.815 0.8 20.815 1.985 21.085 1.985 21.085 2.215 20.115 2.215 20.115 3.155 20.135 3.155 20.135 3.7 19.905 3.7 19.905 3.25 18.005 3.25  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4
