* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I A3:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!((A1 * A2) * A3)
M_i_1_3 net_1_3 A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_0 VSS A3 net_1_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_1 net_1_2 A3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 net_0 A2 net_1_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_1_1 A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_2 VSS A3 net_1_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 net_1_0 A3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 net_0_0 A2 net_1_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_4_3 ZN A2 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_0 VDD A3 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_1 ZN A3 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_4_2 VDD A2 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_4_1 ZN A2 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_2 VDD A3 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_5_3 ZN A3 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_4_0 VDD A2 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_3_3 ZN A1 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_3_2 VDD A1 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_3_1 ZN A1 VDD VNW pmos_5p0 W=1.460000U L=0.500000U
M_i_3_0 VDD A1 ZN VNW pmos_5p0 W=1.460000U L=0.500000U
.ENDS
