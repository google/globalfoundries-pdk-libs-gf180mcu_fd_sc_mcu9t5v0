* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__addh_4 A B CO S VDD VNW VPW VSS
*.PININFO A:I B:I CO:O S:O VDD:P VNW:P VPW:P VSS:G
*.EQN CO=(A * B);S=!((A * B) + !(A + B))
M_i_5_1 net_0_0 A VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4_1 NCO B net_0_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4_0 net_0_1 B NCO VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_5_0 VSS A net_0_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_10_0 net_1 NCO VSS VPW nfet_05v0 W=0.880000U L=0.600000U
M_i_8_0 NS A net_1 VPW nfet_05v0 W=0.880000U L=0.600000U
M_i_9_0 net_1 B NS VPW nfet_05v0 W=0.880000U L=0.600000U
M_i_9_1 NS B net_1 VPW nfet_05v0 W=0.880000U L=0.600000U
M_i_8_1 net_1 A NS VPW nfet_05v0 W=0.880000U L=0.600000U
M_i_10_1 VSS NCO net_1 VPW nfet_05v0 W=0.880000U L=0.600000U
M_i_2_3 CO NCO VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_2 VSS NCO CO VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_1 CO NCO VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_0 VSS NCO CO VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_3 S NS VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_2 VSS NS S VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_1 S NS VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0 VSS NS S VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_7_1 NCO A VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_1 VDD B NCO VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6_0 NCO B VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_7_0 VDD A NCO VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_13_0 NS NCO VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_11_0 net_2_0 A NS VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_12_0 VDD B net_2_0 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_12_1 net_2_1 B VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_11_1 NS A net_2_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_13_1 VDD NCO NS VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_3_3 CO NCO VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_3_2 VDD NCO CO VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_3_1 CO NCO VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_3_0 VDD NCO CO VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_3 S NS VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_2 VDD NS S VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_1 S NS VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_0 VDD NS S VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
