* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I B:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!((A1 * A2) + B)
M_i_1_3 net_0_0 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_3 ZN A1 net_0_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_2 net_0_1 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_2 VSS A2 net_0_1 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_1 net_0_2 A2 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 ZN A1 net_0_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 net_0_3 A1 ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_1_0 VSS A2 net_0_3 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2_3 ZN B VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_2_2 VSS B ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_2_1 ZN B VSS VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_2_0 VSS B ZN VPW nmos_5p0 W=0.920000U L=0.600000U
M_i_4_3 ZN A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_3 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_2 ZN A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_2 net_1 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_1 ZN A2 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_1 net_1 A1 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_3_0 ZN A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_4_0 net_1 A2 ZN VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_3 VDD B net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_2 net_1 B VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_1 VDD B net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5_0 net_1 B VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
