# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.77 1.21 2.695 1.21 2.695 2.115 1.77 2.115  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.626 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.115 1.705 0.97 1.705 0.97 2.595 0.115 2.595  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.925 1.615 3.815 1.615 3.815 2.15 2.925 2.15  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.389 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.045 1.615 4.915 1.615 4.915 2.15 4.045 2.15  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.0102 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.27 0.75 3.28 0.75 3.28 1.06 4.63 1.06 4.63 0.92 4.86 0.92 4.86 1.29 3.05 1.29 3.05 0.98 1.53 0.98 1.53 3.83 1.27 3.83  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 2.52 4.59 4.53 4.59 4.53 3.875 4.76 3.875 4.76 4.59 5.6 4.59 5.6 5.49 2.52 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 3.74 0.45 3.74 0.83 3.51 0.83 3.51 0.45 0.48 0.45 0.48 1.3 0.25 1.3 0.25 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.25 3.55 0.48 3.55 0.48 4.13 2.29 4.13 2.29 3.55 2.52 3.55 2.52 4.36 0.25 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_1
