# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8595 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.21 2.09 1.21 2.09 1.775 4.275 1.775 4.275 2.52 4.045 2.52 4.045 2.005 2.17 2.005 2.17 2.135 1.83 2.135  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8595 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.905 2.18 1.135 2.18 1.135 2.825 2.735 2.825 2.735 2.775 3.31 2.775 4.63 2.775 4.63 2.18 5.295 2.18 5.295 2.71 4.86 2.71 4.86 3.005 3.31 3.005 2.88 3.005 2.88 3.055 0.905 3.055  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.1705 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.91 2.475 9.41 2.475 9.67 2.475 9.67 2.33 10.48 2.33 10.48 2.71 9.41 2.71 7.91 2.71  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.593 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.765 3.235 13.49 3.235 13.72 3.235 13.72 1.72 13.59 1.72 13.59 1.49 12.665 1.49 12.665 0.68 12.895 0.68 12.895 1.21 14.905 1.21 14.905 0.845 15.135 0.845 15.135 1.885 17.145 1.885 17.145 0.845 17.375 0.845 17.375 4.36 17.045 4.36 17.045 2.115 15.185 2.115 15.185 4.36 14.955 4.36 14.955 2.03 13.95 2.03 13.95 3.465 13.49 3.465 12.995 3.465 12.995 4.36 12.765 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.385 4.59 2.385 3.695 2.615 3.695 2.615 4.59 3.31 4.59 5.875 4.59 6.365 4.59 6.365 3.015 6.595 3.015 6.595 4.59 8.685 4.59 8.685 3.865 8.915 3.865 8.915 4.59 11.845 4.59 11.845 4.35 12.075 4.35 12.075 4.59 13.49 4.59 13.785 4.59 13.785 3.695 14.015 3.695 14.015 4.59 15.975 4.59 15.975 3.695 16.205 3.695 16.205 4.59 17.92 4.59 17.92 5.49 13.49 5.49 5.875 5.49 3.31 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 16.255 0.45 16.255 1.655 16.025 1.655 16.025 0.45 14.015 0.45 14.015 0.695 13.785 0.695 13.785 0.45 8.635 0.45 8.635 1.185 8.405 1.185 8.405 0.45 5.875 0.45 5.875 1.185 5.645 1.185 5.645 0.45 2.715 0.45 2.715 1.185 2.485 1.185 2.485 0.45 0.475 0.45 0.475 1.185 0.245 1.185 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 1.72 1.365 1.72 1.365 0.845 1.595 0.845 1.595 2.365 2.38 2.365 2.38 2.235 3.31 2.235 3.31 2.465 2.59 2.465 2.59 2.595 1.365 2.595 1.365 1.95 0.575 1.95 0.575 4.035 0.345 4.035  ;
        POLYGON 3.605 3.695 3.835 3.695 3.835 4.13 5.645 4.13 5.645 3.695 5.875 3.695 5.875 4.36 3.605 4.36  ;
        POLYGON 6.365 0.845 6.595 0.845 6.595 1.72 7.615 1.72 7.615 2.015 9.41 2.015 9.41 2.245 7.615 2.245 7.615 3.22 7.385 3.22 7.385 1.95 6.365 1.95  ;
        POLYGON 4.625 3.235 5.525 3.235 5.525 1.645 4.465 1.645 4.465 1.13 3.55 1.13 3.55 0.9 4.695 0.9 4.695 1.415 5.755 1.415 5.755 2.18 7.055 2.18 7.055 3.45 8.405 3.45 8.405 3.405 11.265 3.405 11.265 2.18 11.495 2.18 11.495 3.635 8.545 3.635 8.545 3.68 6.825 3.68 6.825 2.41 5.755 2.41 5.755 3.465 4.855 3.465 4.855 3.9 4.625 3.9  ;
        POLYGON 9.705 0.68 12.175 0.68 12.175 1.49 11.945 1.49 11.945 0.91 9.935 0.91 9.935 1.655 9.705 1.655  ;
        POLYGON 9.7 3.865 11.725 3.865 11.725 1.95 10.825 1.95 10.825 1.315 11.055 1.315 11.055 1.72 11.955 1.72 11.955 1.93 13.49 1.93 13.49 2.16 11.955 2.16 11.955 4.095 9.7 4.095  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_4
