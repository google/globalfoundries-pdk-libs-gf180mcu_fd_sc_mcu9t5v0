# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__addf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addf_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.04 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.7 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.425 2.33 4.605 2.33 4.605 2.71 3.425 2.71  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.7 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.71 2.15 16.11 2.15 16.11 2.71 14.71 2.71  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.525 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.05 1.92 5.83 1.92 9.135 1.92 13.215 1.92 13.59 1.92 13.59 1.77 13.85 1.77 13.85 2.15 13.215 2.15 9.135 2.15 5.83 2.15 5.05 2.15  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6224 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.165 0.845 17.77 0.845 17.77 2.71 17.395 2.71 17.395 3.685 17.165 3.685  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6224 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 0.845 1.855 0.845 1.855 3.83 1.27 3.83  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.605 4.59 0.605 3.845 0.835 3.845 0.835 4.59 2.645 4.59 2.645 3.845 2.875 3.845 2.875 4.59 5.83 4.59 7.785 4.59 7.785 3.905 8.015 3.905 8.015 4.59 9.035 4.59 10.025 4.59 10.025 3.435 10.255 3.435 10.255 4.59 11.765 4.59 11.765 3.435 11.995 3.435 11.995 4.59 13.115 4.59 15.965 4.59 15.965 3.905 16.195 3.905 16.195 4.59 16.935 4.59 18.185 4.59 18.185 3.845 18.415 3.845 18.415 4.59 19.04 4.59 19.04 5.49 16.935 5.49 13.115 5.49 9.035 5.49 5.83 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.04 -0.45 19.04 0.45 18.735 0.45 18.735 1.165 18.505 1.165 18.505 0.45 16.495 0.45 16.495 1.195 16.265 1.195 16.265 0.45 12.095 0.45 12.095 1.215 11.865 1.215 11.865 0.45 10.255 0.45 10.255 1.215 10.025 1.215 10.025 0.45 8.015 0.45 8.015 1.215 7.785 1.215 7.785 0.45 2.755 0.45 2.755 1.165 2.525 1.165 2.525 0.45 0.515 0.45 0.515 1.165 0.285 1.165 0.285 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.085 1.775 2.965 1.775 2.965 1.37 5.83 1.37 5.83 1.6 3.195 1.6 3.195 2.94 5.545 2.94 5.545 2.875 5.775 2.875 5.775 3.685 5.545 3.685 5.545 3.17 2.965 3.17 2.965 2.115 2.085 2.115  ;
        POLYGON 6.71 2.93 9.035 2.93 9.035 3.74 8.805 3.74 8.805 3.16 6.71 3.16  ;
        POLYGON 6.665 1.315 6.895 1.315 6.895 1.445 8.905 1.445 8.905 1.315 9.135 1.315 9.135 1.675 6.665 1.675  ;
        POLYGON 10.745 2.93 13.115 2.93 13.115 3.74 12.885 3.74 12.885 3.16 10.975 3.16 10.975 3.74 10.745 3.74  ;
        POLYGON 10.745 1.315 10.975 1.315 10.975 1.445 12.985 1.445 12.985 1.315 13.215 1.315 13.215 1.675 10.745 1.675  ;
        POLYGON 6.07 2.47 14.335 2.47 14.335 2.985 16.705 2.985 16.705 1.655 14.05 1.655 14.05 1.37 14.39 1.37 14.39 1.425 16.935 1.425 16.935 3.215 14.105 3.215 14.105 2.7 6.07 2.7  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addf_2
