# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.06 2.39 3.51 2.39 3.51 1.77 3.77 1.77 3.77 1.87 4.79 1.87 4.79 2.39 6.62 2.39 6.62 2.62 4.56 2.62 4.56 2.1 3.77 2.1 3.77 2.62 3.06 2.62  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.87 2.39 1.21 2.39 1.21 2.85 4.07 2.85 4.07 2.33 4.33 2.33 4.33 2.85 6.85 2.85 6.85 2.39 8.81 2.39 8.81 2.62 7.08 2.62 7.08 3.08 0.87 3.08  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.67 2.33 9.955 2.33 9.955 2.85 12.875 2.85 12.875 2.335 13.105 2.335 13.105 2.85 15.24 2.85 15.24 2.39 17.15 2.39 17.15 2.62 15.47 2.62 15.47 3.08 9.67 3.08  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.85 2.39 12.27 2.39 12.27 2 12.33 2 12.33 1.77 13.565 1.77 13.565 2.39 15.01 2.39 15.01 2.62 13.335 2.62 13.335 2 12.73 2 12.73 2.155 12.5 2.155 12.5 2.62 11.85 2.62  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.9601 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.64 3.31 16.655 3.31 16.655 4.36 16.425 4.36 16.425 3.54 14.615 3.54 14.615 4.345 14.385 4.345 14.385 3.54 12.575 3.54 12.575 4.36 12.345 4.36 12.345 3.83 11.91 3.83 11.91 3.54 10.535 3.54 10.535 4.12 10.305 4.12 10.305 3.54 7.145 3.54 7.145 4.36 6.915 4.36 6.915 3.54 2.715 3.54 2.715 4.36 2.485 4.36 2.485 3.54 0.41 3.54 0.41 1.72 1.365 1.72 1.365 1.14 1.595 1.14 1.595 1.72 3.05 1.72 3.05 1.14 4.12 1.14 4.12 1.35 5.845 1.35 5.845 1.14 6.21 1.14 6.21 1.6 8.085 1.6 8.085 1.14 8.315 1.14 8.315 1.83 5.98 1.83 5.98 1.58 3.99 1.58 3.99 1.54 3.28 1.54 3.28 1.95 0.64 1.95  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.77 0.575 3.77 0.575 4.59 4.675 4.59 4.675 3.77 4.905 3.77 4.905 4.59 9.105 4.59 9.105 3.77 9.335 3.77 9.335 4.59 11.325 4.59 11.325 3.77 11.555 3.77 11.555 4.59 13.365 4.59 13.365 3.77 13.595 3.77 13.595 4.59 15.405 4.59 15.405 3.77 15.635 3.77 15.635 4.59 17.445 4.59 17.445 3.77 17.675 3.77 17.675 4.59 17.92 4.59 17.92 5.49 17.675 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 15.635 0.45 15.635 1.49 15.405 1.49 15.405 0.45 11.555 0.45 11.555 1.265 11.325 1.265 11.325 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.68 9.435 0.68 9.435 1.495 11.87 1.495 11.87 1.31 13.365 1.31 13.365 0.68 13.595 0.68 13.595 1.31 14.025 1.31 14.025 1.72 17.445 1.72 17.445 0.68 17.675 0.68 17.675 1.95 13.795 1.95 13.795 1.54 12.1 1.54 12.1 1.725 9.205 1.725 9.205 0.91 7.25 0.91 7.25 0.965 6.91 0.965 6.91 0.91 5.01 0.91 5.01 0.965 4.67 0.965 4.67 0.91 2.77 0.91 2.77 0.965 2.43 0.965 2.43 0.91 0.475 0.91 0.475 1.49 0.245 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_4
