# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 23.52 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.51 2.33 3.995 2.33 3.995 3.27 3.51 3.27  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.144 ;
    PORT
      LAYER METAL1 ;
        POLYGON 18.07 2.89 18.61 2.89 18.61 1.77 18.89 1.77 18.89 3.27 18.07 3.27  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.33 1.53 2.33 1.53 2.735 0.71 2.735  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.77 1.83 2.15 1.83 2.15 2.75 1.77 2.75  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.31 2.33 7.13 2.33 7.13 2.735 6.31 2.735  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6746 ;
    PORT
      LAYER METAL1 ;
        POLYGON 21.895 0.84 22.25 0.84 22.25 4.25 21.895 4.25  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.44 1.595 3.44 1.595 4.59 5.085 4.59 5.085 3.44 5.315 3.44 5.315 4.59 7.175 4.59 7.175 3.94 7.515 3.94 7.515 4.59 9.2 4.59 9.695 4.59 12.03 4.59 12.03 3.44 12.26 3.44 12.26 4.59 13.28 4.59 13.77 4.59 13.77 3.44 13.955 3.44 14 3.44 14 4.59 15.02 4.59 18.07 4.59 18.07 4.48 18.3 4.48 18.3 4.59 20 4.59 20.33 4.59 20.33 3.44 20.56 3.44 20.56 4.59 20.585 4.59 22.915 4.59 22.915 3.44 23.145 3.44 23.145 4.59 23.52 4.59 23.52 5.49 20.585 5.49 20 5.49 15.02 5.49 13.955 5.49 13.28 5.49 9.695 5.49 9.2 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 23.52 -0.45 23.52 0.45 23.275 0.45 23.275 1.16 23.045 1.16 23.045 0.45 21.035 0.45 21.035 1.16 20.805 1.16 20.805 0.45 18.08 0.45 18.08 1.325 17.85 1.325 17.85 0.45 13.36 0.45 13.36 1.325 13.13 1.325 13.13 0.45 7.56 0.45 7.56 1.18 7.33 1.18 7.33 0.45 5.735 0.45 5.735 0.605 5.505 0.605 5.505 0.45 1.595 0.45 1.595 1.14 1.365 1.14 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 2.98 2.545 2.98 2.545 1.6 0.245 1.6 0.245 0.8 0.475 0.8 0.475 1.37 4.99 1.37 4.99 2.735 4.65 2.735 4.65 1.6 2.775 1.6 2.775 3.21 0.575 3.21 0.575 4.25 0.345 4.25  ;
        POLYGON 6.155 2.965 7.36 2.965 7.36 2.1 6.21 2.1 6.21 1.27 6.44 1.27 6.44 1.87 7.59 1.87 7.59 2.505 7.955 2.505 7.955 2.735 7.59 2.735 7.59 3.195 6.155 3.195  ;
        POLYGON 3.125 3.44 3.355 3.44 3.355 4.02 4.625 4.02 4.625 2.98 5.775 2.98 5.775 3.48 8.97 3.48 8.97 3.44 9.2 3.44 9.2 4.25 8.97 4.25 8.97 3.71 5.545 3.71 5.545 3.21 4.855 3.21 4.855 4.25 3.125 4.25  ;
        POLYGON 3.27 0.835 6 0.835 6 0.81 6.9 0.81 6.9 1.41 7.99 1.41 7.99 0.755 9.42 0.755 9.42 1.325 9.19 1.325 9.19 0.985 8.22 0.985 8.22 1.64 6.67 1.64 6.67 1.04 6.105 1.04 6.105 1.065 3.61 1.065 3.61 1.085 3.27 1.085  ;
        POLYGON 8.25 2.52 8.45 2.52 8.45 1.215 8.68 1.215 8.68 2.505 9.695 2.505 9.695 2.735 8.535 2.735 8.535 3.25 8.25 3.25  ;
        POLYGON 11.01 2.98 13.28 2.98 13.28 4.25 13.05 4.25 13.05 3.21 11.24 3.21 11.24 4.25 11.01 4.25  ;
        POLYGON 9.99 2.685 10.31 2.685 10.31 0.985 10.54 0.985 10.54 2.505 13.955 2.505 13.955 2.735 10.535 2.735 10.535 2.915 10.22 2.915 10.22 4.25 9.99 4.25  ;
        POLYGON 11.535 2.045 14.25 2.045 14.25 1.215 14.48 1.215 14.48 3.02 15.02 3.02 15.02 4.25 14.79 4.25 14.79 3.25 14.25 3.25 14.25 2.275 11.535 2.275  ;
        POLYGON 10.835 1.585 13.79 1.585 13.79 0.755 16.5 0.755 16.5 2.79 16.27 2.79 16.27 0.985 15.02 0.985 15.02 2.79 14.79 2.79 14.79 0.985 14.02 0.985 14.02 1.815 11.175 1.815 11.175 1.96 10.835 1.96  ;
        POLYGON 16.73 1.215 17.06 1.215 17.06 3.78 16.73 3.78  ;
        POLYGON 15.39 1.215 16.04 1.215 16.04 4.02 19.77 4.02 19.77 2.525 20 2.525 20 4.25 15.81 4.25 15.81 1.555 15.39 1.555  ;
        POLYGON 17.41 2.45 17.64 2.45 17.64 3.55 19.31 3.55 19.31 1.985 19.99 1.985 19.99 0.8 20.22 0.8 20.22 1.985 20.585 1.985 20.585 2.215 19.54 2.215 19.54 3.78 17.41 3.78  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2
