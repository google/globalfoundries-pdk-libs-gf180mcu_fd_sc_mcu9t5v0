# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 23.52 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.51 2.33 4.525 2.33 4.525 2.71 3.51 2.71  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.71 2.15 15.53 2.15 15.53 2.71 14.71 2.71  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.24 1.575 2.24 1.575 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER METAL1 ;
        POLYGON 19.665 2.875 21.425 2.875 21.655 2.875 21.655 1.655 19.665 1.655 19.665 0.845 19.895 0.845 19.895 1.395 21.43 1.395 21.43 0.815 22.135 0.815 22.135 3.685 21.705 3.685 21.705 3.105 21.425 3.105 19.895 3.105 19.895 3.685 19.665 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.105 4.59 3.105 3.86 3.335 3.86 3.335 4.59 7.345 4.59 7.345 3.905 7.575 3.905 7.575 4.59 9.825 4.59 9.825 3.905 10.055 3.905 10.055 4.59 11.795 4.59 14.205 4.59 14.205 3.915 14.435 3.915 14.435 4.59 16.745 4.59 16.745 3.155 16.975 3.155 16.975 4.59 17.47 4.59 18.645 4.59 18.645 3.875 18.875 3.875 18.875 4.59 20.685 4.59 20.685 3.875 20.915 3.875 20.915 4.59 21.425 4.59 22.725 4.59 22.725 3.875 22.955 3.875 22.955 4.59 23.52 4.59 23.52 5.49 21.425 5.49 17.47 5.49 11.795 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 23.52 -0.45 23.52 0.45 23.255 0.45 23.255 1.165 23.025 1.165 23.025 0.45 21.015 0.45 21.015 1.165 20.785 1.165 20.785 0.45 18.775 0.45 18.775 1.165 18.545 1.165 18.545 0.45 16.755 0.45 16.755 1.425 16.525 1.425 16.525 0.45 7.755 0.45 7.755 1.425 7.525 1.425 7.525 0.45 3.455 0.45 3.455 1.425 3.225 1.425 3.225 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 1.685 0.245 1.685 0.245 1.315 0.475 1.315 0.475 1.455 2.035 1.455 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 3.28 2.94 4.63 2.94 4.63 3.205 4.29 3.205 4.29 3.17 3.05 3.17 3.05 1.87 4.345 1.87 4.345 1.315 4.575 1.315 4.575 2.1 3.28 2.1  ;
        POLYGON 5.365 1.315 5.795 1.315 5.795 1.83 8.29 1.83 8.29 2.06 5.595 2.06 5.595 3.26 5.365 3.26  ;
        POLYGON 6.63 2.515 9.825 2.515 9.825 1.315 10.055 1.315 10.055 2.515 11.355 2.515 11.355 3.215 11.125 3.215 11.125 2.745 8.815 2.745 8.815 3.215 8.585 3.215 8.585 2.745 6.63 2.745  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 3.4 3.705 3.4 3.705 3.49 5.895 3.49 5.895 3.445 11.795 3.445 11.795 4.315 11.565 4.315 11.565 3.675 6.035 3.675 6.035 4.36 5.805 4.36 5.805 3.72 3.52 3.72 3.52 3.63 2.615 3.63 2.615 3.685 2.385 3.685  ;
        POLYGON 13.485 2.875 14.105 2.875 14.105 1.545 12.245 1.545 12.245 1.205 14.335 1.205 14.335 2.995 15.79 2.995 15.79 3.225 13.485 3.225  ;
        POLYGON 11.125 1.315 11.355 1.315 11.355 1.775 12.375 1.775 12.375 3.455 16.285 3.455 16.285 2.48 17.47 2.48 17.47 2.71 16.515 2.71 16.515 3.685 12.145 3.685 12.145 2.005 11.125 2.005  ;
        POLYGON 16.085 1.775 17.825 1.775 17.825 1.315 18.055 1.315 18.055 1.96 21.425 1.96 21.425 2.32 17.995 2.32 17.995 3.695 17.765 3.695 17.765 2.115 16.085 2.115  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4
