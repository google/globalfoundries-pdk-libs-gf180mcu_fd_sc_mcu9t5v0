# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.8 1.71 11.73 1.71 11.73 2.15 9.8 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.825 2.325 1.055 2.325 1.055 2.895 3.51 2.895 3.51 2.33 3.77 2.33 3.77 2.38 4.33 2.38 4.33 2.895 6.745 2.895 6.745 2.38 8.81 2.38 8.81 2.61 6.975 2.61 6.975 3.125 0.825 3.125  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.556 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.94 1.77 6.515 1.77 6.515 2.665 6.285 2.665 6.285 2.15 4.07 2.15 4.07 2 3.28 2 3.28 2.61 2.94 2.61  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.734 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.325 2.65 11.96 2.65 11.96 1.48 1.365 1.48 1.365 0.68 1.595 0.68 1.595 1.25 3.605 1.25 3.605 0.68 3.835 0.68 3.835 1.25 5.845 1.25 5.845 0.68 6.075 0.68 6.075 1.25 8.085 1.25 8.085 0.68 8.315 0.68 8.315 1.25 10.325 1.25 10.325 0.68 10.555 0.68 10.555 1.25 12.565 1.25 12.565 0.68 12.795 0.68 12.795 1.48 12.19 1.48 12.19 3.09 12.695 3.09 12.695 3.9 11.91 3.9 11.91 2.88 10.555 2.88 10.555 3.9 10.325 3.9  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 2.385 4.59 2.385 3.825 2.615 3.825 2.615 4.59 6.865 4.59 6.865 3.815 7.095 3.815 7.095 4.59 13.815 4.59 14.56 4.59 14.56 5.49 13.815 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 13.915 0.45 13.915 1.02 13.685 1.02 13.685 0.45 11.675 0.45 11.675 1.02 11.445 1.02 11.445 0.45 9.435 0.45 9.435 1.02 9.205 1.02 9.205 0.45 7.195 0.45 7.195 1.02 6.965 1.02 6.965 0.45 4.955 0.45 4.955 1.02 4.725 1.02 4.725 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.02 0.245 1.02 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 3.11 0.475 3.11 0.475 3.355 7.605 3.355 7.605 4.13 11.345 4.13 11.345 3.11 11.575 3.11 11.575 4.13 13.585 4.13 13.585 3.11 13.815 3.11 13.815 4.36 7.375 4.36 7.375 3.585 4.855 3.585 4.855 4.165 4.625 4.165 4.625 3.585 0.475 3.585 0.475 3.92 0.245 3.92  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__nor3_4
