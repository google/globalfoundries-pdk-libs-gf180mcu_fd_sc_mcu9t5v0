# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__addh_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.3 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.1 2.215 1.33 2.215 1.33 2.63 3.93 2.63 3.93 2.285 6.45 2.285 6.45 2.63 7.85 2.63 7.85 2.27 9.86 2.27 9.86 2.5 8.08 2.5 8.08 2.86 1.1 2.86  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.3 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.77 1.825 6.91 1.825 6.91 2.17 7.62 2.17 7.62 2.4 6.68 2.4 6.68 2.055 3.05 2.055 3.05 2.4 1.77 2.4  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.5505 ;
    PORT
      LAYER METAL1 ;
        POLYGON 12.47 1.365 15.15 1.365 15.15 1.595 12.805 1.595 12.805 2.985 15.1 2.985 15.1 3.215 12.47 3.215  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.6603 ;
    PORT
      LAYER METAL1 ;
        POLYGON 16.95 2.96 18.59 2.96 19.075 2.96 19.075 1.79 16.95 1.79 16.95 0.695 17.335 0.695 17.335 1.43 19.345 1.43 19.345 0.695 19.575 0.695 19.575 1.79 19.435 1.79 19.435 4.36 19.205 4.36 19.205 3.32 18.59 3.32 17.235 3.32 17.235 4.36 16.95 4.36  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 2.335 4.59 2.335 3.55 2.565 3.55 2.565 4.59 4.425 4.59 4.425 3.55 4.655 3.55 4.655 4.59 7.915 4.59 7.915 4.01 8.145 4.01 8.145 4.59 11.275 4.59 11.275 4.01 11.505 4.01 11.505 4.59 13.695 4.59 13.695 4.01 13.925 4.01 13.925 4.59 15.885 4.59 15.885 3.55 16.115 3.55 16.115 4.59 18.125 4.59 18.125 3.55 18.355 3.55 18.355 4.59 18.59 4.59 20.335 4.59 20.335 3.55 20.565 3.55 20.565 4.59 21.28 4.59 21.28 5.49 18.59 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.695 0.45 20.695 1.2 20.465 1.2 20.465 0.45 18.455 0.45 18.455 1.2 18.225 1.2 18.225 0.45 16.215 0.45 16.215 1.2 15.985 1.2 15.985 0.675 11.735 0.675 11.735 1.125 11.505 1.125 11.505 0.45 4.655 0.45 4.655 1.595 4.425 1.595 4.425 0.45 0.475 0.45 0.475 1.2 0.245 1.2 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 5.67 0.845 10.49 0.845 10.49 1.075 5.67 1.075  ;
        POLYGON 0.87 3.09 10.09 3.09 10.09 2.27 12.23 2.27 12.23 2.5 10.32 2.5 10.32 3.32 3.635 3.32 3.635 4.36 3.405 4.36 3.405 3.32 1.545 3.32 1.545 4.36 1.315 4.36 1.315 3.32 0.64 3.32 0.64 1.365 2.385 1.365 2.385 0.695 2.615 0.695 2.615 1.595 0.87 1.595  ;
        POLYGON 5.725 3.55 15.38 3.55 15.38 1.135 12.195 1.135 12.195 1.585 6.79 1.585 6.79 1.355 11.965 1.355 11.965 0.905 15.61 0.905 15.61 2.215 18.59 2.215 18.59 2.555 15.61 2.555 15.61 3.78 10.385 3.78 10.385 4.36 10.155 4.36 10.155 3.78 5.955 3.78 5.955 4.36 5.725 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_4
