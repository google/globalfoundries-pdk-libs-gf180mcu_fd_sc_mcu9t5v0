# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.6 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.43 2.33 4.33 2.33 4.33 2.71 3.43 2.71  ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.33 1.705 2.33 1.705 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER METAL1 ;
        POLYGON 15.71 2.89 17.555 2.89 17.785 2.89 17.785 1.64 15.71 1.64 15.71 1.37 18.29 1.37 18.29 3.23 17.555 3.23 15.71 3.23  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.495 4.59 1.495 3.425 1.725 3.425 1.725 4.59 2.165 4.59 3.435 4.59 3.435 3.515 3.665 3.515 3.665 4.59 6.3 4.59 7.535 4.59 7.535 3.045 7.765 3.045 7.765 4.59 9.265 4.59 12.805 4.59 12.805 4.345 13.035 4.345 13.035 4.59 14.745 4.59 14.745 4.345 14.975 4.345 14.975 4.59 16.785 4.59 16.785 4.345 17.015 4.345 17.015 4.59 18.75 4.59 18.825 4.59 18.825 4.345 19.055 4.345 19.055 4.59 19.6 4.59 19.6 5.49 18.75 5.49 9.265 5.49 6.3 5.49 2.165 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 19.6 -0.45 19.6 0.45 19.355 0.45 19.355 1.165 19.125 1.165 19.125 0.45 17.17 0.45 17.17 0.64 16.83 0.64 16.83 0.45 14.93 0.45 14.93 0.64 14.59 0.64 14.59 0.45 13.09 0.45 13.09 0.64 12.75 0.64 12.75 0.45 7.985 0.45 7.985 0.625 7.755 0.625 7.755 0.45 3.565 0.45 3.565 1.145 3.335 1.145 3.335 0.45 1.725 0.45 1.725 1.225 1.495 1.225 1.495 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.475 2.94 1.935 2.94 1.935 2.005 0.375 2.005 0.375 1.315 0.605 1.315 0.605 1.775 2.165 1.775 2.165 3.17 0.705 3.17 0.705 3.75 0.475 3.75  ;
        POLYGON 4.555 2.875 4.56 2.875 4.56 1.375 4.455 1.375 4.455 1.035 4.79 1.035 4.79 3.685 4.555 3.685  ;
        POLYGON 2.515 1.315 2.845 1.315 2.845 2.985 4.125 2.985 4.125 4.03 6.3 4.03 6.3 4.26 3.895 4.26 3.895 3.215 2.515 3.215  ;
        POLYGON 5.575 1.035 5.805 1.035 5.805 2.01 8.355 2.01 8.355 1.9 8.585 1.9 8.585 2.24 5.805 2.24 5.805 3.685 5.575 3.685  ;
        POLYGON 7.04 2.47 9.035 2.47 9.035 1.315 9.265 1.315 9.265 3.685 9.03 3.685 9.03 2.7 7.04 2.7  ;
        POLYGON 6.2 0.855 9.42 0.855 9.42 0.68 11.395 0.68 11.395 2.755 11.165 2.755 11.165 1.085 6.54 1.085 6.54 1.78 6.2 1.78  ;
        POLYGON 10.155 1.315 10.385 1.315 10.385 2.985 11.625 2.985 11.625 2.47 13.53 2.47 13.53 2.7 11.855 2.7 11.855 3.215 10.385 3.215 10.385 3.685 10.155 3.685  ;
        POLYGON 12.31 1.92 13.87 1.92 13.87 1.37 14.21 1.37 14.21 1.87 17.555 1.87 17.555 2.21 14.055 2.21 14.055 3.215 13.825 3.215 13.825 2.15 12.31 2.15  ;
        POLYGON 11.73 3.5 18.52 3.5 18.52 1.14 11.915 1.14 11.915 1.49 11.685 1.49 11.685 0.68 11.915 0.68 11.915 0.91 18.75 0.91 18.75 3.73 11.73 3.73  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_4
