# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai22_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 10.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.28 2.27 6.62 2.27 6.62 2.71 6.28 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.35 2.27 5.69 2.27 5.69 2.94 6.87 2.94 6.87 2.215 8.755 2.215 8.755 3.17 5.35 3.17  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.75 2.27 2.09 2.27 2.09 2.71 1.75 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.87 2.27 1.21 2.27 1.21 2.94 2.39 2.94 2.39 2.27 4.33 2.27 4.33 3.17 0.87 3.17  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.7335 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.535 3.4 8.985 3.4 8.985 1.985 5.845 1.985 5.845 1.14 6.075 1.14 6.075 1.755 7.99 1.755 7.99 1.14 8.315 1.14 8.315 1.755 9.215 1.755 9.215 3.63 7.145 3.63 7.145 4.36 6.915 4.36 6.915 3.63 2.765 3.63 2.765 4.36 2.535 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.86 0.575 3.86 0.575 4.59 4.625 4.59 4.625 3.86 4.855 3.86 4.855 4.59 9.105 4.59 9.105 3.86 9.335 3.86 9.335 4.59 9.435 4.59 10.08 4.59 10.08 5.49 9.435 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 10.08 -0.45 10.08 0.45 3.835 0.45 3.835 1.055 3.605 1.055 3.605 0.45 1.595 0.45 1.595 1.525 1.365 1.525 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.715 0.475 0.715 0.475 1.755 2.485 1.755 2.485 1.285 4.725 1.285 4.725 0.68 9.435 0.68 9.435 1.525 9.205 1.525 9.205 0.91 7.195 0.91 7.195 1.525 6.965 1.525 6.965 0.91 4.955 0.91 4.955 1.985 0.245 1.985  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai22_2
