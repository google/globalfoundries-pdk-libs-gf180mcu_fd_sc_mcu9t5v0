# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 21.28 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.83 1.96 4.63 1.96 4.63 1.77 4.89 1.77 4.89 2.19 3.83 2.19  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.655 2.165 14.86 2.165 14.86 2.71 13.655 2.71  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.235 1.575 2.235 1.575 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.12 0.845 19.45 0.845 19.45 3.685 19.12 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.305 4.59 3.305 3.58 3.535 3.58 3.535 4.59 7.305 4.59 7.305 3.11 7.535 3.11 7.535 4.59 9.365 4.59 9.365 3.11 9.595 3.11 9.595 4.59 11.435 4.59 13.745 4.59 13.745 3.97 13.975 3.97 13.975 4.59 16.345 4.59 16.345 3.21 16.575 3.21 16.575 4.59 17.07 4.59 18.1 4.59 18.1 3.875 18.33 3.875 18.33 4.59 18.77 4.59 20.14 4.59 20.14 3.875 20.37 3.875 20.37 4.59 21.28 4.59 21.28 5.49 18.77 5.49 17.07 5.49 11.435 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 21.28 -0.45 21.28 0.45 20.57 0.45 20.57 1.165 20.34 1.165 20.34 0.45 18.33 0.45 18.33 1.165 18.1 1.165 18.1 0.45 16.475 0.45 16.475 1.42 16.245 1.42 16.245 0.45 7.635 0.45 7.635 1.325 7.405 1.325 7.405 0.45 3.49 0.45 3.49 1.27 3.15 1.27 3.15 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.9 0.575 2.9 0.575 2.94 1.805 2.94 1.805 2.005 0.245 2.005 0.245 1.315 0.475 1.315 0.475 1.775 2.035 1.775 2.035 3.17 0.575 3.17 0.575 3.71 0.345 3.71  ;
        POLYGON 3.6 2.42 4.555 2.42 4.555 3.75 4.325 3.75 4.325 2.65 3.37 2.65 3.37 1.5 3.715 1.5 3.715 1.32 4.325 1.32 4.325 1.21 4.555 1.21 4.555 1.55 3.94 1.55 3.94 1.73 3.6 1.73  ;
        POLYGON 5.445 1.215 5.675 1.215 5.675 1.73 8.13 1.73 8.13 1.96 5.675 1.96 5.675 3.75 5.445 3.75  ;
        POLYGON 6.81 2.19 9.365 2.19 9.365 1.215 9.595 1.215 9.595 2.19 10.995 2.19 10.995 3.685 10.765 3.685 10.765 2.42 8.555 2.42 8.555 3.75 8.325 3.75 8.325 2.42 6.81 2.42  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 2.985 3.995 2.985 3.995 4.095 6.845 4.095 6.845 2.65 7.995 2.65 7.995 3.98 8.905 3.98 8.905 2.65 10.055 2.65 10.055 3.975 11.435 3.975 11.435 4.315 9.825 4.315 9.825 2.88 9.135 2.88 9.135 4.21 7.765 4.21 7.765 2.88 7.075 2.88 7.075 4.325 3.765 4.325 3.765 3.215 2.385 3.215  ;
        POLYGON 13.255 2.94 15.275 2.94 15.275 3.28 13.025 3.28 13.025 1.5 11.785 1.5 11.785 1.16 13.875 1.16 13.875 1.5 13.255 1.5  ;
        POLYGON 10.665 1.215 10.895 1.215 10.895 1.73 12.015 1.73 12.015 3.51 15.885 3.51 15.885 2.535 17.07 2.535 17.07 2.765 16.115 2.765 16.115 3.74 11.785 3.74 11.785 1.96 10.665 1.96  ;
        POLYGON 15.625 1.775 17.365 1.775 17.365 1.315 17.595 1.315 17.595 1.775 18.77 1.775 18.77 2.115 17.595 2.115 17.595 3.75 17.365 3.75 17.365 2.115 15.625 2.115  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2
