* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__and2_4 A1 A2 Z VDD VNW VPW VSS
*.PININFO A1:I A2:I Z:O VDD:P VNW:P VPW:P VSS:G
*.EQN Z=(A1 * A2)
M_i_3_1 net_0_1 A2 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_1 Z_neg A1 net_0_1 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2_0 net_0_0 A1 Z_neg VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3_0 VSS A2 net_0_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_3 Z Z_neg VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_2 VSS Z_neg Z VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_1 Z Z_neg VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0_0 VSS Z_neg Z VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_5_1 Z_neg A2 VDD VNW pfet_05v0 W=1.640000U L=0.500000U
M_i_4_1 VDD A1 Z_neg VNW pfet_05v0 W=1.640000U L=0.500000U
M_i_4_0 Z_neg A1 VDD VNW pfet_05v0 W=1.640000U L=0.500000U
M_i_5_0 VDD A2 Z_neg VNW pfet_05v0 W=1.640000U L=0.500000U
M_i_1_3 Z Z_neg VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_2 VDD Z_neg Z VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_1 Z Z_neg VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_1_0 VDD Z_neg Z VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
