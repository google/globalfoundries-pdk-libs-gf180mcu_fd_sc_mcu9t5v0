# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.692 ;
    PORT
      LAYER METAL1 ;
        POLYGON 7.99 1.77 8.46 1.77 8.46 2.71 7.99 2.71  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6224 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.62 0.68 6.85 0.68 6.85 1.21 7.13 1.21 7.13 2.71 7 2.71 7 3.75 6.77 3.75 6.77 1.49 6.62 1.49  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.37 4.59 1.37 3.4 1.6 3.4 1.6 4.59 5.75 4.59 5.75 4.35 5.98 4.35 5.98 4.59 7.79 4.59 7.79 3.4 8.02 3.4 8.02 4.59 9.09 4.59 9.52 4.59 9.52 5.49 9.09 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 7.97 0.45 7.97 1.49 7.74 1.49 7.74 0.45 5.73 0.45 5.73 1.02 5.5 1.02 5.5 0.45 1.65 0.45 1.65 1.02 1.42 1.02 1.42 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.35 2.94 1.86 2.94 1.86 1.49 0.3 1.49 0.3 0.68 0.53 0.68 0.53 1.26 2.09 1.26 2.09 2.47 3.625 2.47 3.625 3.17 0.58 3.17 0.58 4.21 0.35 4.21  ;
        POLYGON 2.54 0.68 5.265 0.68 5.265 1.25 6.39 1.25 6.39 2.11 6.16 2.11 6.16 1.48 5.035 1.48 5.035 1.085 3.43 1.085 3.43 2.01 4.15 2.01 4.15 3.9 3.92 3.9 3.92 2.24 3.2 2.24 3.2 1.49 2.54 1.49  ;
        POLYGON 2.9 3.4 3.13 3.4 3.13 4.13 4.585 4.13 4.585 1.78 3.66 1.78 3.66 1.315 3.89 1.315 3.89 1.55 4.815 1.55 4.815 1.99 5.93 1.99 5.93 2.465 6.475 2.465 6.475 2.695 5.7 2.695 5.7 2.22 4.96 2.22 4.96 4.36 2.9 4.36  ;
        POLYGON 5.24 2.45 5.47 2.45 5.47 2.925 6.395 2.925 6.395 3.98 7.33 3.98 7.33 2.94 8.86 2.94 8.86 0.68 9.09 0.68 9.09 4.21 8.81 4.21 8.81 3.17 7.56 3.17 7.56 4.21 6.165 4.21 6.165 3.155 5.24 3.155  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_2
