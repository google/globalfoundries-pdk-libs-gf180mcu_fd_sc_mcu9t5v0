# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.698 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 2.015 0.97 2.015 0.97 2.71 0.15 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.849 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.505 1.77 8.81 1.77 8.81 2.71 8.505 2.71  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.3728 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.61 1.14 4.84 1.14 4.84 1.77 4.89 1.77 4.89 3.9 4.61 3.9  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.48 1.495 3.48 1.495 4.59 5.68 4.59 5.68 3.86 5.91 3.86 5.91 4.59 6.795 4.59 7.585 4.59 7.585 3.48 7.815 3.48 7.815 4.59 9.33 4.59 9.52 4.59 9.52 5.49 9.33 5.49 6.795 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 7.815 0.45 7.815 1.48 7.585 1.48 7.585 0.45 5.96 0.45 5.96 1.165 5.73 1.165 5.73 0.45 1.84 0.45 1.84 1.48 1.61 1.48 1.61 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 3.02 2.105 3.02 2.105 2.245 1.2 2.245 1.2 1.82 1.095 1.82 1.095 1.425 0.19 1.425 0.19 1.195 1.325 1.195 1.325 1.625 1.43 1.625 1.43 2.015 2.335 2.015 2.335 3.02 3.06 3.02 3.06 3.25 0.475 3.25 0.475 4.29 0.245 4.29  ;
        POLYGON 2.675 1.195 3.355 1.195 3.355 0.68 5.3 0.68 5.3 1.395 6.465 1.395 6.465 1.14 6.695 1.14 6.695 1.625 5.375 1.625 5.375 2.17 5.145 2.17 5.145 1.565 5.07 1.565 5.07 0.91 3.585 0.91 3.585 3.82 3.355 3.82 3.355 1.425 2.675 1.425  ;
        POLYGON 2.335 3.48 2.565 3.48 2.565 4.13 3.85 4.13 3.85 1.14 4.08 1.14 4.08 4.13 5.12 4.13 5.12 2.43 5.415 2.43 5.415 3.4 6.795 3.4 6.795 4.29 6.565 4.29 6.565 3.63 5.35 3.63 5.35 4.36 2.335 4.36  ;
        POLYGON 7.09 2.015 8.045 2.015 8.045 1.195 9.33 1.195 9.33 1.425 8.275 1.425 8.275 3.15 9.175 3.15 9.175 4.29 8.945 4.29 8.945 3.38 8.045 3.38 8.045 2.245 7.09 2.245  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_1
