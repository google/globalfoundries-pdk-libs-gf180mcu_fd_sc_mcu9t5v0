* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__icgtp_2 CLK E TE Q VDD VNW VPW VSS
*.PININFO CLK:I E:I TE:I Q:O VDD:P VNW:P VPW:P VSS:G
M_MU19 net50 TE VSS VPW nfet_05v0 W=0.700000U L=0.600000U
M_MU20 VSS E net50 VPW nfet_05v0 W=0.700000U L=0.600000U
M_MI82 net50 NCK net53 VPW nfet_05v0 W=0.700000U L=0.600000U
M_MI91 net53 CK net033 VPW nfet_05v0 W=0.700000U L=0.600000U
M_MI92 net033 QD VSS VPW nfet_05v0 W=0.700000U L=0.600000U
M_MI80_M_u2 VSS net53 QD VPW nfet_05v0 W=0.700000U L=0.600000U
M_MU82_M_u2 VSS NCK CK VPW nfet_05v0 W=0.700000U L=0.600000U
M_MU81_M_u2 NCK CLK VSS VPW nfet_05v0 W=0.700000U L=0.600000U
M_MI85_M_u3 XI85-net6 CLK d3 VPW nfet_05v0 W=1.000000U L=0.600000U
M_MI85_M_u4 VSS QD XI85-net6 VPW nfet_05v0 W=1.000000U L=0.600000U
M_MU75_M_u2 Q d3 VSS VPW nfet_05v0 W=1.000000U L=0.600000U
M_MU75_M_u2_22 Q d3 VSS VPW nfet_05v0 W=1.000000U L=0.600000U
M_MI81 VDD TE net58 VNW pfet_05v0 W=1.380000U L=0.500000U
M_MU17 net58 E net61 VNW pfet_05v0 W=1.380000U L=0.500000U
M_MU16 net61 CK net53 VNW pfet_05v0 W=1.380000U L=0.500000U
M_MI90 net53 NCK net062 VNW pfet_05v0 W=1.380000U L=0.500000U
M_MI88 net062 QD VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_MI80_M_u3 VDD net53 QD VNW pfet_05v0 W=1.380000U L=0.500000U
M_MU82_M_u3 CK NCK VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_MU81_M_u3 VDD CLK NCK VNW pfet_05v0 W=1.380000U L=0.500000U
M_MI85_M_u1 d3 CLK VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_MI85_M_u2 VDD QD d3 VNW pfet_05v0 W=1.830000U L=0.500000U
M_MU75_M_u3 Q d3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_MU75_M_u3_3 Q d3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
