# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai32_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai32_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.32 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 2.27 3.26 2.27 3.26 2.71 2.92 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 2.27 2.46 2.27 2.46 1.81 4.63 1.81 4.63 1.77 4.89 1.77 4.89 2.27 5.45 2.27 5.45 2.5 4.63 2.5 4.63 2.04 2.69 2.04 2.69 2.5 1.94 2.5  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.94 5.68 2.94 5.68 2.27 6.57 2.27 6.57 2.5 5.91 2.5 5.91 3.17 0.71 3.17  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.515 2.215 8.81 2.215 8.81 2.71 8.515 2.71  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.43 2.215 7.735 2.215 7.735 2.94 10.765 2.94 10.765 2.215 10.995 2.215 10.995 3.17 7.43 3.17  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.655 3.415 11.225 3.415 11.225 1.985 7.99 1.985 7.99 1.14 8.315 1.14 8.315 1.755 10.325 1.755 10.325 1.14 10.555 1.14 10.555 1.755 11.455 1.755 11.455 3.645 9.385 3.645 9.385 4.34 9.155 4.34 9.155 3.645 3.885 3.645 3.885 4.355 3.655 4.355  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.875 0.575 3.875 0.575 4.59 6.865 4.59 6.865 3.875 7.095 3.875 7.095 4.59 11.345 4.59 11.345 3.875 11.575 3.875 11.575 4.59 11.915 4.59 12.32 4.59 12.32 5.49 11.915 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 12.32 -0.45 12.32 0.45 6.075 0.45 6.075 1.095 5.845 1.095 5.845 0.45 3.835 0.45 3.835 1.095 3.605 1.095 3.605 0.45 1.595 0.45 1.595 1.095 1.365 1.095 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.755 0.475 0.755 0.475 1.335 2.485 1.335 2.485 0.755 2.715 0.755 2.715 1.335 4.37 1.335 4.37 1.31 4.725 1.31 4.725 0.73 5.16 0.73 5.16 1.335 6.965 1.335 6.965 0.68 11.915 0.68 11.915 1.565 11.685 1.565 11.685 0.91 9.435 0.91 9.435 1.525 9.205 1.525 9.205 0.91 7.195 0.91 7.195 1.565 5.055 1.565 5.055 1.54 4.475 1.54 4.475 1.565 0.245 1.565  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai32_2
