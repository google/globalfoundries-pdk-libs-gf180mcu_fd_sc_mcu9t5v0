# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 28 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.656 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.44 2.27 7.83 2.27 7.83 2.65 0.44 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 14.568 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.325 2.96 16.98 2.96 17.805 2.96 17.805 2.04 10.325 2.04 10.325 0.68 10.555 0.68 10.555 1.72 12.565 1.72 12.565 0.68 12.795 0.68 12.795 1.72 14.805 1.72 14.805 0.68 15.035 0.68 15.035 1.72 17.045 1.72 17.045 0.68 17.305 0.68 17.305 1.72 19.285 1.72 19.285 0.68 19.515 0.68 19.515 1.72 21.525 1.72 21.525 0.68 21.755 0.68 21.755 1.72 23.765 1.72 23.765 0.68 23.995 0.68 23.995 1.72 26.005 1.72 26.005 0.68 26.235 0.68 26.235 1.985 18.555 1.985 18.555 2.96 26.065 2.96 26.135 2.96 26.135 4.36 26.065 4.36 25.905 4.36 25.905 3.32 23.895 3.32 23.895 4.36 23.665 4.36 23.665 3.32 21.655 3.32 21.655 4.36 21.425 4.36 21.425 3.32 19.415 3.32 19.415 4.36 19.185 4.36 19.185 3.32 17.175 3.32 17.175 4.36 16.98 4.36 16.945 4.36 16.945 3.32 14.935 3.32 14.935 4.36 14.705 4.36 14.705 3.32 12.695 3.32 12.695 4.36 12.465 4.36 12.465 3.32 10.555 3.32 10.555 4.36 10.325 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.55 11.575 3.55 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 15.825 4.59 15.825 3.55 16.055 3.55 16.055 4.59 16.98 4.59 18.065 4.59 18.065 3.55 18.295 3.55 18.295 4.59 20.305 4.59 20.305 3.55 20.535 3.55 20.535 4.59 22.545 4.59 22.545 3.55 22.775 3.55 22.775 4.59 24.785 4.59 24.785 3.55 25.015 3.55 25.015 4.59 26.065 4.59 27.025 4.59 27.025 3.55 27.255 3.55 27.255 4.59 28 4.59 28 5.49 26.065 5.49 16.98 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 28 -0.45 28 0.45 27.355 0.45 27.355 1.49 27.125 1.49 27.125 0.45 25.115 0.45 25.115 1.49 24.885 1.49 24.885 0.45 22.875 0.45 22.875 1.49 22.645 1.49 22.645 0.45 20.635 0.45 20.635 1.49 20.405 1.49 20.405 0.45 18.395 0.45 18.395 1.49 18.165 1.49 18.165 0.45 16.155 0.45 16.155 1.49 15.925 1.49 15.925 0.45 13.915 0.45 13.915 1.49 13.685 1.49 13.685 0.45 11.675 0.45 11.675 1.49 11.445 1.49 11.445 0.45 9.435 0.45 9.435 1.49 9.205 1.49 9.205 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.88 8.06 2.88 8.06 2.04 1.365 2.04 1.365 0.68 1.595 0.68 1.595 1.72 3.605 1.72 3.605 0.68 3.835 0.68 3.835 1.72 5.845 1.72 5.845 0.68 6.075 0.68 6.075 1.72 8.085 1.72 8.085 0.68 8.425 0.68 8.425 2.27 16.98 2.27 16.98 2.63 8.425 2.63 8.425 4.36 8.06 4.36 8.06 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
        POLYGON 18.785 2.215 26.065 2.215 26.065 2.555 18.785 2.555  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_16
