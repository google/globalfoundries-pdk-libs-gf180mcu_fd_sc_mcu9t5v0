# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 26.88 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 1.77 4.33 1.77 4.33 2.29 3.51 2.29  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.123 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.43 1.77 21.69 1.77 21.69 2.015 21.935 2.015 21.935 2.355 21.69 2.355 21.69 2.71 21.43 2.71  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.77 0.97 1.77 0.97 2.3 0.15 2.3  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.75 1.77 20.04 1.77 20.04 2.71 19.75 2.71  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 1.77 2.09 1.77 2.09 2.345 1.27 2.345  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.31 2.33 7.13 2.33 7.13 2.71 6.31 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 25.145 0.79 25.61 0.79 25.61 2.71 25.375 2.71 25.375 4.08 25.145 4.08  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.415 4.59 1.415 3.27 1.645 3.27 1.645 4.59 5.085 4.59 5.085 3.44 5.315 3.44 5.315 4.59 7.19 4.59 7.19 4.125 7.53 4.125 7.53 4.59 9.215 4.59 9.655 4.59 9.695 4.59 12.21 4.59 12.21 4.565 12.55 4.565 12.55 4.59 15.35 4.59 15.35 4.565 15.69 4.565 15.69 4.59 17.31 4.59 19.395 4.59 19.395 3.91 19.625 3.91 19.625 4.59 21.665 4.59 21.665 4.3 21.895 4.3 21.895 4.59 23.375 4.59 23.725 4.59 23.725 3.27 23.955 3.27 23.955 4.59 24.835 4.59 26.165 4.59 26.165 3.27 26.395 3.27 26.395 4.59 26.88 4.59 26.88 5.49 24.835 5.49 23.375 5.49 17.31 5.49 9.695 5.49 9.655 5.49 9.215 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 26.88 -0.45 26.88 0.45 26.635 0.45 26.635 1.6 26.405 1.6 26.405 0.45 24.395 0.45 24.395 1.6 24.165 1.6 24.165 0.45 21.31 0.45 21.31 1.08 20.97 1.08 20.97 0.45 13.775 0.45 13.775 1.48 13.545 1.48 13.545 0.45 7.775 0.45 7.775 1.08 7.545 1.08 7.545 0.45 5.735 0.45 5.735 1.08 5.505 1.08 5.505 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.395 2.575 2.595 2.575 2.595 1.54 0.245 1.54 0.245 0.79 0.475 0.79 0.475 1.31 2.825 1.31 2.825 2.52 4.605 2.52 4.605 2.015 4.835 2.015 4.835 2.75 2.745 2.75 2.745 2.805 0.625 2.805 0.625 4.08 0.395 4.08  ;
        POLYGON 6.225 3.095 7.36 3.095 7.36 2 6.425 2 6.425 1.17 6.655 1.17 6.655 1.77 8.215 1.77 8.215 2.11 7.59 2.11 7.59 3.435 6.225 3.435  ;
        POLYGON 3.325 2.98 5.775 2.98 5.775 3.665 8.985 3.665 8.985 3.085 9.215 3.085 9.215 3.895 5.545 3.895 5.545 3.21 3.555 3.21 3.555 4.08 3.325 4.08  ;
        POLYGON 8.265 2.335 8.665 2.335 8.665 1.17 8.895 1.17 8.895 2.225 9.655 2.225 9.655 2.565 8.495 2.565 8.495 3.435 8.265 3.435  ;
        POLYGON 3.325 0.79 3.555 0.79 3.555 1.31 5.965 1.31 5.965 0.71 7.115 0.71 7.115 1.31 8.205 1.31 8.205 0.71 9.695 0.71 9.695 1.48 9.465 1.48 9.465 0.94 8.435 0.94 8.435 1.54 6.885 1.54 6.885 0.94 6.195 0.94 6.195 1.54 3.325 1.54  ;
        POLYGON 11.025 3.27 13.675 3.27 13.675 3.61 11.025 3.61  ;
        POLYGON 10.005 2.74 10.585 2.74 10.585 1.37 10.815 1.37 10.815 2.74 14.535 2.74 14.535 3.08 14.305 3.08 14.305 2.97 10.235 2.97 10.235 3.93 10.005 3.93  ;
        POLYGON 14.165 3.535 15.905 3.535 15.905 2.51 12.005 2.51 12.005 2.17 15.905 2.17 15.905 1.37 16.135 1.37 16.135 3.645 16.585 3.645 16.585 3.065 16.815 3.065 16.815 3.875 14.165 3.875  ;
        POLYGON 10.53 4.105 17.31 4.105 17.31 4.335 10.53 4.335  ;
        POLYGON 11.165 1.71 15.445 1.71 15.445 0.68 18.835 0.68 18.835 2.355 18.605 2.355 18.605 1.02 15.675 1.02 15.675 1.94 11.395 1.94 11.395 2.355 11.165 2.355  ;
        POLYGON 18.145 1.37 18.375 1.37 18.375 2.585 19.065 2.585 19.065 1.025 19.295 1.025 19.295 1.31 20.63 1.31 20.63 3.27 20.645 3.27 20.645 3.61 20.4 3.61 20.4 1.54 19.295 1.54 19.295 2.815 18.855 2.815 18.855 3.305 18.625 3.305 18.625 2.815 18.145 2.815  ;
        POLYGON 17.025 1.37 17.255 1.37 17.255 2.74 17.835 2.74 17.835 3.535 19.035 3.535 19.035 3.45 20.085 3.45 20.085 3.84 23.145 3.84 23.145 2.415 23.375 2.415 23.375 4.07 19.855 4.07 19.855 3.68 19.215 3.68 19.215 3.765 17.605 3.765 17.605 2.97 17.025 2.97  ;
        POLYGON 20.86 1.31 23.445 1.31 23.445 0.845 23.675 0.845 23.675 1.965 24.835 1.965 24.835 2.355 24.605 2.355 24.605 2.195 23.445 2.195 23.445 1.54 22.915 1.54 22.915 3.61 22.685 3.61 22.685 1.54 21.2 1.54 21.2 2.3 20.86 2.3  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2
