# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__and4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.28 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.115 2.15 0.97 2.15 0.97 2.71 0.115 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.2 2.15 2.09 2.15 2.09 2.71 1.2 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.32 2.29 3.21 2.29 3.21 2.71 2.32 2.71  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.432 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.44 2.33 4.33 2.33 4.33 2.71 3.44 2.71  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.19 0.845 6.1 0.845 6.1 3.685 5.58 3.685 5.58 1.725 5.19 1.725  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.3 4.59 0.3 3.875 0.53 3.875 0.53 4.59 2.34 4.59 2.34 4.345 2.57 4.345 2.57 4.59 4.38 4.59 4.38 3.875 4.61 3.875 4.61 4.59 5.23 4.59 6.6 4.59 6.6 3.875 6.83 3.875 6.83 4.59 7.28 4.59 7.28 5.49 5.23 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 7.28 -0.45 7.28 0.45 6.85 0.45 6.85 1.165 6.62 1.165 6.62 0.45 4.61 0.45 4.61 0.695 4.38 0.695 4.38 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.32 3.415 4.56 3.415 4.56 1.6 0.245 1.6 0.245 1.37 4.79 1.37 4.79 2.38 5.23 2.38 5.23 2.72 4.79 2.72 4.79 3.645 3.59 3.645 3.59 4.235 3.36 4.235 3.36 3.765 1.32 3.765  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and4_2
