# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 14.56 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 16.236 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.63 2.27 6.14 2.27 6.14 2.65 0.63 2.65  ;
        POLYGON 7.66 2.27 13.17 2.27 13.17 2.65 7.66 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.0852 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.365 3.09 6.37 3.09 6.37 1.745 1.365 1.745 1.365 0.945 1.595 0.945 1.595 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 5.845 1.515 5.845 0.945 6.075 0.945 6.075 1.515 8.085 1.515 8.085 0.945 8.315 0.945 8.315 1.515 10.325 1.515 10.325 0.945 10.555 0.945 10.555 1.515 12.565 1.515 12.565 0.945 12.795 0.945 12.795 1.745 7.12 1.745 7.12 3.09 12.695 3.09 12.695 4.36 12.465 4.36 12.465 3.32 10.455 3.32 10.455 4.36 10.225 4.36 10.225 3.32 8.215 3.32 8.215 4.36 7.985 4.36 7.985 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.55 9.335 3.55 9.335 4.59 11.345 4.59 11.345 3.55 11.575 3.55 11.575 4.59 13.585 4.59 13.585 3.55 13.815 3.55 13.815 4.59 14.56 4.59 14.56 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 14.56 -0.45 14.56 0.45 13.915 0.45 13.915 1.285 13.685 1.285 13.685 0.45 11.675 0.45 11.675 1.285 11.445 1.285 11.445 0.45 9.435 0.45 9.435 1.285 9.205 1.285 9.205 0.45 7.195 0.45 7.195 1.285 6.965 1.285 6.965 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_12
