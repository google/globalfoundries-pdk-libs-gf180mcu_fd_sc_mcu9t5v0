# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nand4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.96 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.51 2.215 3.875 2.215 3.875 2.71 3.51 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.865 2.215 3.095 2.215 3.095 2.94 4.235 2.94 4.235 2.215 6.015 2.215 6.015 2.71 4.465 2.71 4.465 3.17 2.865 3.17  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.755 7.035 1.755 7.035 2.555 6.805 2.555 6.805 1.985 2.09 1.985 2.09 2.555 1.83 2.555  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.864 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.825 2.215 1.27 2.215 1.27 1.77 1.53 1.77 1.53 3.31 2.235 3.31 2.235 3.4 4.695 3.4 4.695 2.94 7.825 2.94 7.825 2.215 8.055 2.215 8.055 3.17 4.925 3.17 4.925 3.63 2.05 3.63 2.05 3.54 1.3 3.54 1.3 2.555 0.825 2.555  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.8096 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.475 3.77 1.865 3.77 1.865 3.86 5.065 3.86 5.065 3.815 6.365 3.815 6.365 3.4 8.635 3.4 8.635 4.36 8.405 4.36 8.405 3.63 6.595 3.63 6.595 4.045 5.205 4.045 5.205 4.09 1.68 4.09 1.68 4 0.475 4 0.475 4.36 0.15 4.36 0.15 1.755 0.81 1.755 0.81 0.68 4.555 0.68 4.555 1.49 4.325 1.49 4.325 0.91 1.04 0.91 1.04 1.985 0.475 1.985  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 4.23 1.495 4.23 1.495 4.59 3.305 4.59 3.305 4.32 3.535 4.32 3.535 4.59 5.345 4.59 5.345 4.275 5.575 4.275 5.575 4.59 7.385 4.59 7.385 3.86 7.615 3.86 7.615 4.59 8.96 4.59 8.96 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 8.96 -0.45 8.96 0.45 8.635 0.45 8.635 1.49 8.405 1.49 8.405 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand4_2
