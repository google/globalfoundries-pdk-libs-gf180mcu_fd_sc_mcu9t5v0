# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__xor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.88 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.89 1.77 2.42 1.77 2.42 1.41 4.455 1.41 4.455 2.21 4.225 2.21 4.225 1.64 2.65 1.64 2.65 2.155 1.89 2.155  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.925 1.87 1.155 1.87 1.155 2.845 3.335 2.845 5.245 2.845 5.245 1.87 5.475 1.87 5.475 3.075 3.335 3.075 1.53 3.075 1.53 3.27 0.925 3.27  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER METAL1 ;
        POLYGON 7.99 2.33 8.335 2.33 8.335 2.48 9.74 2.48 10.525 2.48 10.525 1.87 10.755 1.87 10.755 2.71 9.74 2.71 7.99 2.71  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.105 2.89 11.775 2.89 12.005 2.89 12.005 1.155 10.03 1.155 10.03 0.895 10.37 0.895 10.37 0.925 12.235 0.925 12.235 3.27 11.775 3.27 11.335 3.27 11.335 3.7 11.105 3.7  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 2.385 4.59 2.385 3.305 2.615 3.305 2.615 4.59 3.335 4.59 6.11 4.59 8.685 4.59 8.685 2.965 8.915 2.965 8.915 4.59 9.74 4.59 12.635 4.59 12.88 4.59 12.88 5.49 12.635 5.49 9.74 5.49 6.11 5.49 3.335 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 12.88 -0.45 12.88 0.45 12.355 0.45 12.355 0.695 12.125 0.695 12.125 0.45 9.015 0.45 9.015 1.18 8.785 1.18 8.785 0.45 6.775 0.45 6.775 1.18 6.545 1.18 6.545 0.45 6.055 0.45 6.055 1.18 5.825 1.18 5.825 0.45 2.715 0.45 2.715 1.18 2.485 1.18 2.485 0.45 0.475 0.45 0.475 1.18 0.245 1.18 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 1.41 1.365 1.41 1.365 0.84 1.615 0.84 1.615 2.385 3.105 2.385 3.105 1.87 3.335 1.87 3.335 2.615 1.385 2.615 1.385 1.64 0.575 1.64 0.575 3.645 0.345 3.645  ;
        POLYGON 3.785 3.305 4.015 3.305 4.015 3.83 6.11 3.83 6.11 4.115 3.785 4.115  ;
        POLYGON 6.63 2.44 7.53 2.44 7.53 1.89 7.665 1.89 7.665 1.14 7.895 1.14 7.895 1.87 9.74 1.87 9.74 2.155 9.4 2.155 9.4 2.1 7.76 2.1 7.76 2.67 6.86 2.67 6.86 3.775 6.63 3.775  ;
        POLYGON 4.75 3.36 5.705 3.36 5.705 1.64 4.685 1.64 4.685 1.125 3.73 1.125 3.73 0.895 4.915 0.895 4.915 1.41 7.205 1.41 7.205 0.68 8.555 0.68 8.555 1.41 11.775 1.41 11.775 2.21 11.545 2.21 11.545 1.64 8.325 1.64 8.325 0.91 7.435 0.91 7.435 1.62 7.3 1.62 7.3 2.21 7.07 2.21 7.07 1.64 5.935 1.64 5.935 3.59 4.75 3.59  ;
        POLYGON 10.085 3.305 10.315 3.305 10.315 4.005 12.405 4.005 12.405 3.425 12.635 3.425 12.635 4.235 10.085 4.235  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor3_1
