# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.706 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.805 1.77 1.53 1.77 1.53 2.215 1.975 2.215 1.975 2.555 0.805 2.555  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.1012 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.785 3.09 4.745 3.09 5.75 3.09 5.75 1.675 3.785 1.675 3.785 0.875 4.015 0.875 4.015 1.445 5.75 1.445 5.75 0.875 6.255 0.875 6.255 1.875 6.155 1.875 6.155 4.36 5.925 4.36 5.925 3.32 4.745 3.32 4.015 3.32 4.015 4.36 3.785 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.745 4.59 4.805 4.59 4.805 3.55 5.035 3.55 5.035 4.59 7.045 4.59 7.045 3.55 7.275 3.55 7.275 4.59 7.84 4.59 7.84 5.49 4.745 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 7.375 0.45 7.375 1.215 7.145 1.215 7.145 0.45 5.135 0.45 5.135 1.215 4.905 1.215 4.905 0.45 2.895 0.45 2.895 1.215 2.665 1.215 2.665 0.45 0.475 0.45 0.475 1.215 0.245 1.215 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 3.09 2.205 3.09 2.205 1.16 1.31 1.16 1.31 0.93 2.435 0.93 2.435 2.215 4.745 2.215 4.745 2.555 2.435 2.555 2.435 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_4
