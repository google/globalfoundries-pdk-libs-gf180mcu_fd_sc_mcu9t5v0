# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__clkinv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkinv_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.059 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 2.215 1.83 2.215 1.83 1.77 2.09 1.77 2.09 2.215 2.325 2.215 2.325 2.71 0.685 2.71  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.6406 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.09 3.51 3.09 3.51 1.44 1.365 1.44 1.365 0.68 1.595 0.68 1.595 1.21 3.605 1.21 3.605 0.68 3.835 0.68 3.835 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.48 4.59 4.48 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 2.715 0.45 2.715 0.98 2.485 0.98 2.485 0.45 0.475 0.45 0.475 1.02 0.245 1.02 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__clkinv_3
