# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dlyd_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlyd_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 18.48 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.66 1.77 1 1.77 1 2.595 0.66 2.595  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.825 ;
    PORT
      LAYER METAL1 ;
        POLYGON 14.695 2.89 16.13 2.89 16.36 2.89 16.36 1.9 14.645 1.9 14.645 0.68 14.875 0.68 14.875 1.67 16.885 1.67 16.885 0.68 17.115 0.68 17.115 1.9 16.59 1.9 16.59 2.89 16.965 2.89 16.965 4.36 16.735 4.36 16.735 3.12 16.13 3.12 14.97 3.12 14.97 4.36 14.695 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.275 4.59 1.275 3.93 1.505 3.93 1.505 4.59 4.395 4.59 4.745 4.59 4.745 3.93 4.975 3.93 4.975 4.59 8.395 4.59 8.745 4.59 8.745 3.93 8.975 3.93 8.975 4.59 12.395 4.59 12.745 4.59 12.745 3.93 12.975 3.93 12.975 4.59 15.715 4.59 15.715 3.88 15.945 3.88 15.945 4.59 16.13 4.59 17.905 4.59 17.905 3.88 18.135 3.88 18.135 4.59 18.48 4.59 18.48 5.49 16.13 5.49 12.395 5.49 8.395 5.49 4.395 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 18.48 -0.45 18.48 0.45 18.235 0.45 18.235 1.44 18.005 1.44 18.005 0.45 15.995 0.45 15.995 1.44 15.765 1.44 15.765 0.45 13.075 0.45 13.075 0.695 12.845 0.695 12.845 0.45 9.075 0.45 9.075 0.965 8.845 0.965 8.845 0.45 5.075 0.45 5.075 0.97 4.845 0.97 4.845 0.45 1.605 0.45 1.605 0.97 1.375 0.97 1.375 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.43 2.825 1.32 2.825 1.32 2.805 1.95 2.805 1.95 1.895 2.29 1.895 2.29 3.035 1.415 3.035 1.415 3.055 0.485 3.055 0.485 4.27 0.2 4.27 0.2 0.685 0.54 0.685 0.54 0.915 0.43 0.915  ;
        POLYGON 1.51 3.265 2.52 3.265 2.52 1.635 1.51 1.635 1.51 1.405 4.395 1.405 4.395 2.65 4.165 2.65 4.165 1.635 2.75 1.635 2.75 3.495 1.51 3.495  ;
        POLYGON 4.745 1.35 5.075 1.35 5.075 1.895 6.29 1.895 6.29 2.595 5.95 2.595 5.95 2.125 4.975 2.125 4.975 3.55 4.745 3.55  ;
        POLYGON 5.565 2.825 6.52 2.825 6.52 1.635 5.51 1.635 5.51 1.405 8.395 1.405 8.395 2.65 8.165 2.65 8.165 1.635 6.75 1.635 6.75 3.055 5.795 3.055 5.795 3.55 5.565 3.55  ;
        POLYGON 8.745 1.345 9.075 1.345 9.075 1.895 10.29 1.895 10.29 2.595 9.95 2.595 9.95 2.125 8.975 2.125 8.975 3.55 8.745 3.55  ;
        POLYGON 9.565 2.825 10.52 2.825 10.52 1.63 9.51 1.63 9.51 1.4 10.75 1.4 10.75 1.84 12.395 1.84 12.395 2.65 12.165 2.65 12.165 2.07 10.75 2.07 10.75 3.055 9.795 3.055 9.795 3.55 9.565 3.55  ;
        POLYGON 12.745 1.075 13.075 1.075 13.075 2.13 16.13 2.13 16.13 2.36 12.975 2.36 12.975 3.55 12.745 3.55  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlyd_4
