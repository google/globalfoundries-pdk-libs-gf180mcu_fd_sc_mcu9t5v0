# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__latsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.32 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.21 2.09 1.21 2.09 2.335 1.83 2.335  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.925 1.995 1.155 1.995 1.155 2.565 2.95 2.565 2.95 1.77 3.21 1.77 3.21 2.05 3.465 2.05 3.465 3.09 4.08 3.09 4.08 3.32 3.235 3.32 3.235 2.795 0.925 2.795  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.87 1.77 7.155 1.77 7.155 2.71 6.87 2.71  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.575 0.68 11.05 0.68 11.05 2.15 10.805 2.15 10.805 4.2 10.575 4.2  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.415 4.59 1.415 3.665 1.645 3.665 1.645 4.59 3.005 4.59 5.115 4.59 5.115 3.55 5.345 3.55 5.345 4.59 7.335 4.59 7.335 3.55 7.565 3.55 7.565 4.59 9.555 4.59 9.555 3.86 9.785 3.86 9.785 4.59 10.225 4.59 11.595 4.59 11.595 3.55 11.825 3.55 11.825 4.59 12.32 4.59 12.32 5.49 10.225 5.49 3.005 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 12.32 -0.45 12.32 0.45 12.075 0.45 12.075 1.49 11.845 1.49 11.845 0.45 9.835 0.45 9.835 1.305 9.605 1.305 9.605 0.45 5.695 0.45 5.695 1.02 5.465 1.02 5.465 0.45 1.595 0.45 1.595 1.02 1.365 1.02 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 3.025 3.005 3.025 3.005 3.365 0.625 3.365 0.625 4.36 0.245 4.36  ;
        POLYGON 3.355 3.55 3.585 3.55 3.585 4.13 4.31 4.13 4.31 1.765 3.505 1.765 3.505 0.68 3.735 0.68 3.735 1.535 5.965 1.535 5.965 2.335 5.735 2.335 5.735 1.765 4.54 1.765 4.54 4.36 3.355 4.36  ;
        POLYGON 5.025 1.995 5.255 1.995 5.255 2.94 8.975 2.94 8.975 2.225 7.605 2.225 7.605 0.68 7.835 0.68 7.835 1.995 9.205 1.995 9.205 3.17 6.545 3.17 6.545 4.2 6.315 4.2 6.315 3.17 5.025 3.17  ;
        POLYGON 8.535 3.4 9.995 3.4 9.995 1.765 8.485 1.765 8.485 0.68 8.715 0.68 8.715 1.535 10.225 1.535 10.225 3.63 8.765 3.63 8.765 4.21 8.535 4.21  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latsnq_2
