# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__mux2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.4 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 1.77 6.57 1.77 6.57 2.15 5.75 2.15  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 1.77 3.255 1.77 3.255 2.71 2.95 2.71  ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.005 1.775 4.235 1.775 4.235 2.47 6.87 2.47 6.87 1.77 7.315 1.77 7.315 2.71 4.005 2.71  ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7295 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 0.68 1.595 0.68 1.595 4.36 1.27 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 5.115 4.59 6.645 4.59 6.645 3.55 6.875 3.55 6.875 4.59 7.995 4.59 8.4 4.59 8.4 5.49 7.995 5.49 5.115 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.4 -0.45 8.4 0.45 6.875 0.45 6.875 1.02 6.645 1.02 6.645 0.45 2.715 0.45 2.715 1.02 2.485 1.02 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.175 2.94 5.115 2.94 5.115 4.36 4.885 4.36 4.885 3.17 1.945 3.17 1.945 1.31 4.445 1.31 4.445 0.68 4.675 0.68 4.675 1.54 2.175 1.54  ;
        POLYGON 4.83 1.83 5.29 1.83 5.29 1.31 7.765 1.31 7.765 0.68 7.995 0.68 7.995 4.36 7.665 4.36 7.665 1.54 5.52 1.54 5.52 2.06 4.83 2.06  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux2_2
