# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 16.8 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 2.33 4.33 2.33 4.33 2.71 3.45 2.71  ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.235 1.57 2.235 1.57 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.71 1.315 15.055 1.315 15.055 3.215 14.71 3.215  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.035 4.59 3.305 4.59 3.305 3.61 3.535 3.61 3.535 4.59 6.17 4.59 7.405 4.59 7.405 3.14 7.635 3.14 7.635 4.59 9.195 4.59 12.545 4.59 12.545 3.905 12.775 3.905 12.775 4.59 15.515 4.59 15.845 4.59 15.845 3.875 16.075 3.875 16.075 4.59 16.8 4.59 16.8 5.49 15.515 5.49 9.195 5.49 6.17 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 16.8 -0.45 16.8 0.45 16.175 0.45 16.175 1.165 15.945 1.165 15.945 0.45 12.995 0.45 12.995 0.625 12.765 0.625 12.765 0.45 7.855 0.45 7.855 0.625 7.625 0.625 7.625 0.45 3.435 0.45 3.435 1.13 3.205 1.13 3.205 0.45 1.595 0.45 1.595 1.225 1.365 1.225 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.94 1.805 2.94 1.805 1.74 0.245 1.74 0.245 1.315 0.475 1.315 0.475 1.51 2.035 1.51 2.035 3.17 0.575 3.17 0.575 3.75 0.345 3.75  ;
        POLYGON 4.425 2.97 4.56 2.97 4.56 1.36 4.325 1.36 4.325 1.02 4.79 1.02 4.79 3.78 4.425 3.78  ;
        POLYGON 2.385 1.315 2.715 1.315 2.715 2.99 3.995 2.99 3.995 4.125 6.17 4.125 6.17 4.355 3.765 4.355 3.765 3.22 2.385 3.22  ;
        POLYGON 5.445 1.02 5.675 1.02 5.675 2.05 8.285 2.05 8.285 1.94 8.515 1.94 8.515 2.28 5.675 2.28 5.675 3.78 5.445 3.78  ;
        POLYGON 6.965 2.51 8.965 2.51 8.965 1.315 9.195 1.315 9.195 3.78 8.965 3.78 8.965 2.85 6.965 2.85  ;
        POLYGON 6.125 0.855 9.35 0.855 9.35 0.68 10.775 0.68 10.775 2.3 11.25 2.3 11.25 2.53 10.545 2.53 10.545 1.085 6.355 1.085 6.355 1.82 6.125 1.82  ;
        POLYGON 10.085 1.315 10.315 1.315 10.315 2.76 13.41 2.76 13.41 2.99 10.315 2.99 10.315 3.78 10.085 3.78  ;
        POLYGON 12.05 2.23 14.105 2.23 14.105 1.315 14.48 1.315 14.48 2.455 14.155 2.455 14.155 3.215 13.925 3.215 13.925 2.46 12.05 2.46  ;
        POLYGON 11.47 3.445 15.285 3.445 15.285 1.085 11.655 1.085 11.655 1.225 11.425 1.225 11.425 0.855 15.515 0.855 15.515 3.675 11.47 3.675  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_1
