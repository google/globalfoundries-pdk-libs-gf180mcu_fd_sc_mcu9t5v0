* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(((A1 + A2) + A3) * ((B1 + B2) + B3))
M_i_5 net_0 B3 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_4 VSS B2 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_3 net_0 B1 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_0 ZN A1 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_1 net_0 A2 ZN VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_2 ZN A3 net_0 VPW nfet_05v0 W=1.320000U L=0.600000U
M_i_11 net_4 B3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_10 net_3 B2 net_4 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_9 ZN B1 net_3 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_6 net_1 A1 ZN VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_7 net_2 A2 net_1 VNW pfet_05v0 W=1.830000U L=0.500000U
M_i_8 VDD A3 net_2 VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
