# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__xnor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xnor3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.88 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.995 1.815 2.225 1.815 2.225 2.33 3.44 2.33 3.67 2.33 3.67 1.87 4.51 1.87 4.51 2.1 3.9 2.1 3.9 2.71 3.44 2.71 1.995 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.317 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.87 1.77 1.53 1.77 1.53 2.94 3.44 2.94 5.245 2.94 5.245 1.815 5.475 1.815 5.475 3.17 3.44 3.17 1.3 3.17 1.3 2.15 0.87 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.09 1.87 8.97 1.87 8.97 2.33 9.54 2.33 9.77 2.33 9.77 1.87 10.71 1.87 10.71 2.1 10 2.1 10 2.71 9.54 2.71 8.74 2.71 8.74 2.1 8.09 2.1  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9125 ;
    PORT
      LAYER METAL1 ;
        POLYGON 9.985 3.49 11.685 3.49 11.685 3.415 11.73 3.415 11.96 3.415 11.96 1.59 10.95 1.59 10.95 1.21 12.19 1.21 12.19 3.645 11.855 3.645 11.855 3.72 11.73 3.72 10.215 3.72 10.215 4.36 9.985 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.55 2.665 3.55 2.665 4.59 3.44 4.59 6.055 4.59 6.545 4.59 6.545 3.855 6.775 3.855 6.775 4.59 8.815 4.59 8.815 3.875 9.045 3.875 9.045 4.59 11.73 4.59 12.025 4.59 12.025 3.875 12.255 3.875 12.255 4.59 12.41 4.59 12.88 4.59 12.88 5.49 12.41 5.49 11.73 5.49 6.055 5.49 3.44 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 12.88 -0.45 12.88 0.45 8.815 0.45 8.815 1.08 8.585 1.08 8.585 0.45 6.055 0.45 6.055 1.08 5.825 1.08 5.825 0.45 2.715 0.45 2.715 1.08 2.485 1.08 2.485 0.45 0.475 0.45 0.475 1.08 0.245 1.08 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.345 1.31 1.365 1.31 1.365 0.74 1.595 0.74 1.595 1.31 2.685 1.31 2.685 1.87 3.44 1.87 3.44 2.1 2.455 2.1 2.455 1.54 0.575 1.54 0.575 3.89 0.345 3.89  ;
        POLYGON 3.785 3.55 4.015 3.55 4.015 4.13 5.825 4.13 5.825 3.855 6.055 3.855 6.055 4.36 3.785 4.36  ;
        POLYGON 6.545 1.04 6.775 1.04 6.775 1.41 9.54 1.41 9.54 2.1 9.2 2.1 9.2 1.64 7.795 1.64 7.795 3.64 7.565 3.64 7.565 1.64 6.545 1.64  ;
        POLYGON 5.955 3.395 7.235 3.395 7.235 3.87 8.355 3.87 8.355 3.03 11.285 3.03 11.285 1.87 11.73 1.87 11.73 2.1 11.515 2.1 11.515 3.26 8.585 3.26 8.585 4.1 7.005 4.1 7.005 3.625 5.775 3.625 5.775 3.63 5.035 3.63 5.035 3.89 4.805 3.89 4.805 3.4 5.725 3.4 5.725 1.54 3.785 1.54 3.785 0.74 4.015 0.74 4.015 1.31 5.955 1.31 5.955 1.87 7.27 1.87 7.27 2.1 5.955 2.1  ;
        POLYGON 9.885 0.74 12.41 0.74 12.41 0.97 10.115 0.97 10.115 1.55 9.885 1.55  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xnor3_1
