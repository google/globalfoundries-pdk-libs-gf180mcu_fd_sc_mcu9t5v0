* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__bufz_16 EN I Z VDD VNW VPW VSS
*.PININFO EN:I I:I Z:O VDD:P VNW:P VPW:P VSS:G
*.EQN Z=I
M_mn VSS EN NEN VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn8 NI_N NEN VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn21 NI_P EN NI_N VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn17 NI_N I VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn17_9 VSS I NI_N VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn17_10 NI_N I VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn17_9_17 VSS I NI_N VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn17_34 NI_N I VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn17_9_41 VSS I NI_N VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn17_10_30 NI_N I VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn17_9_17_61 VSS I NI_N VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_1_25_34 Z NI_N VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_49_88 VSS NI_N Z VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_1_33 Z NI_N VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_99 VSS NI_N Z VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_1_25 Z NI_N VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_49 VSS NI_N Z VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_1 Z NI_N VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3 VSS NI_N Z VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_1_25_34_75 Z NI_N VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_49_88_82 VSS NI_N Z VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_1_33_198 Z NI_N VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_99_125 VSS NI_N Z VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_1_25_137 Z NI_N VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_49_181 VSS NI_N Z VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_1_65 Z NI_N VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_mn3_118 VSS NI_N Z VPW nfet_05v0 W=1.320000U L=0.600000U
M_mp VDD EN NEN VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp7 NI_P EN VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp22 NI_N NEN NI_P VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp14 NI_P I VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp14_10 VDD I NI_P VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp14_11 NI_P I VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp14_10_8 VDD I NI_P VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp14_7 NI_P I VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp14_10_32 VDD I NI_P VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp14_11_55 NI_P I VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp14_10_8_20 VDD I NI_P VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_12_57_75 Z NI_P VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_56_111 VDD NI_P Z VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_12_106 Z NI_P VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_58 VDD NI_P Z VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_12_57 Z NI_P VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_56 VDD NI_P Z VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_12 Z NI_P VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4 VDD NI_P Z VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_12_57_75_85 Z NI_P VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_56_111_134 VDD NI_P Z VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_12_106_111 Z NI_P VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_58_95 VDD NI_P Z VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_12_57_97 Z NI_P VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_56_133 VDD NI_P Z VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_12_126 Z NI_P VDD VNW pfet_05v0 W=1.800000U L=0.500000U
M_mp4_153 VDD NI_P Z VNW pfet_05v0 W=1.800000U L=0.500000U
.ENDS
