# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__inv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__inv_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.58 2.27 2.33 2.27 2.33 2.65 0.58 2.65  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 3.12 3.335 3.12 3.335 1.89 1.365 1.89 1.365 0.68 1.595 0.68 1.595 1.66 3.605 1.66 3.605 0.68 3.835 0.68 3.835 4.36 3.505 4.36 3.505 3.35 1.595 3.35 1.595 4.36 1.365 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.58 2.615 3.58 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 5.6 4.59 5.6 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 4.955 0.45 4.955 1.43 4.725 1.43 4.725 0.45 2.715 0.45 2.715 1.43 2.485 1.43 2.485 0.45 0.475 0.45 0.475 1.43 0.245 1.43 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__inv_4
