# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nor2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.934 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 2.27 2.14 2.27 2.14 2.71 1.8 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.934 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.875 2.215 1.105 2.215 1.105 2.94 3.51 2.94 3.51 1.77 3.77 1.77 3.77 2.27 3.95 2.27 3.95 3.17 0.875 3.17  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9999 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.485 3.55 4.18 3.55 4.18 1.72 4.07 1.72 4.07 1.49 1.365 1.49 1.365 0.68 1.595 0.68 1.595 1.16 3.605 1.16 3.605 0.68 3.835 0.68 3.835 1.21 4.41 1.21 4.41 3.78 2.715 3.78 2.715 4.36 2.485 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 4.675 4.59 4.675 3.55 4.905 3.55 4.905 4.59 5.6 4.59 5.6 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 4.955 0.45 4.955 1.4 4.725 1.4 4.725 0.45 2.715 0.45 2.715 0.93 2.485 0.93 2.485 0.45 0.475 0.45 0.475 1.4 0.245 1.4 0.245 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nor2_2
