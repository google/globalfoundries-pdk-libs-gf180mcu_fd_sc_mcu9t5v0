# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.035 2.215 4.33 2.215 4.33 2.71 4.035 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.95 2.27 3.31 2.27 3.31 2.94 6.285 2.94 6.285 2.215 6.515 2.215 6.515 3.17 2.95 3.17  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.229 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.65 2.27 1.07 2.27 1.07 2.65 0.65 2.65  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.3628 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.365 3.4 6.745 3.4 6.745 1.95 3.605 1.95 3.605 1.14 3.835 1.14 3.835 1.72 5.19 1.72 5.19 1.14 6.075 1.14 6.075 1.72 6.975 1.72 6.975 3.63 4.905 3.63 4.905 4.36 4.675 4.36 4.675 3.63 1.595 3.63 1.595 4.32 1.365 4.32  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.665 0.575 3.665 0.575 4.59 2.385 4.59 2.385 3.86 2.615 3.86 2.615 4.59 6.865 4.59 6.865 3.86 7.095 3.86 7.095 4.59 7.195 4.59 7.84 4.59 7.84 5.49 7.195 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 1.595 0.45 1.595 1.49 1.365 1.49 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.68 0.475 0.68 0.475 1.72 2.485 1.72 2.485 0.68 7.195 0.68 7.195 1.49 6.965 1.49 6.965 0.91 4.955 0.91 4.955 1.49 4.725 1.49 4.725 0.91 2.715 0.91 2.715 1.95 0.245 1.95  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_2
