# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__mux4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__mux4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.36 BY 5.04 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.71 1.21 14.97 1.21 14.97 2.555 14.71 2.555  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.35 1.77 11.61 1.77 11.61 2.71 11.35 2.71  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8535 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.07 1.77 4.375 1.77 4.375 2.71 4.07 2.71  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 1.67 3.21 1.67 3.21 1.9 2.65 1.9 2.65 2.995 2.39 2.995  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.675 1.77 8.105 1.77 8.81 1.77 8.81 3.195 8.405 3.195 8.405 2.155 8.105 2.155 7.675 2.155  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0032 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.75 2.33 6.025 2.33 6.025 1.59 5.75 1.59 5.75 1.21 6.255 1.21 6.255 3.175 5.75 3.175  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.44 0.525 3.44 0.525 4.59 1.595 4.59 4.725 4.59 4.725 3.865 4.955 3.865 4.955 4.59 7.035 4.59 8.105 4.59 10.935 4.59 10.935 3.44 11.165 3.44 11.165 4.59 13.305 4.59 15.015 4.59 15.015 3.44 15.245 3.44 15.245 4.59 16.665 4.59 17.36 4.59 17.36 5.49 16.665 5.49 13.305 5.49 8.105 5.49 7.035 5.49 1.595 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.36 -0.45 17.36 0.45 15.545 0.45 15.545 1.43 15.315 1.43 15.315 0.45 11.065 0.45 11.065 1.43 10.835 1.43 10.835 0.45 4.955 0.45 4.955 1.43 4.725 1.43 4.725 0.45 0.475 0.45 0.475 1.43 0.245 1.43 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 1.09 1.595 1.09 1.595 4.17 1.365 4.17  ;
        POLYGON 3.605 1.09 3.835 1.09 3.835 3.355 3.915 3.355 3.915 3.695 3.605 3.695  ;
        POLYGON 2.16 3.225 2.895 3.225 2.895 3.94 4.265 3.94 4.265 3.405 6.755 3.405 6.755 1.155 6.985 1.155 6.985 3.36 7.035 3.36 7.035 4.17 6.805 4.17 6.805 3.635 4.495 3.635 4.495 4.17 2.665 4.17 2.665 3.455 1.93 3.455 1.93 1.145 2.77 1.145 2.77 1.375 2.16 1.375  ;
        POLYGON 5.29 0.695 8.105 0.695 8.105 1.345 7.875 1.345 7.875 0.925 7.445 0.925 7.445 2.385 8.055 2.385 8.055 4.17 7.825 4.17 7.825 2.615 7.215 2.615 7.215 0.925 5.52 0.925 5.52 1.79 5.575 1.79 5.575 2.13 5.29 2.13  ;
        POLYGON 9.5 1.09 10.145 1.09 10.145 3.695 9.915 3.695 9.915 2.315 9.5 2.315  ;
        POLYGON 11.955 1.09 12.185 1.09 12.185 3.695 11.955 3.695  ;
        POLYGON 8.845 3.425 9.04 3.425 9.04 1.43 8.995 1.43 8.995 1.09 9.27 1.09 9.27 4.005 10.475 4.005 10.475 2.98 11.625 2.98 11.625 3.94 12.975 3.94 12.975 1.09 13.305 1.09 13.305 4.17 11.395 4.17 11.395 3.21 10.705 3.21 10.705 4.235 8.845 4.235  ;
        POLYGON 13.675 1.145 14.48 1.145 14.48 1.375 13.905 1.375 13.905 3.245 14.225 3.245 14.225 4.25 13.995 4.25 13.995 3.475 13.675 3.475  ;
        POLYGON 14.135 2.215 14.365 2.215 14.365 2.785 16.435 2.785 16.435 1.09 16.665 1.09 16.665 3.015 16.265 3.015 16.265 4.17 16.035 4.17 16.035 3.015 14.135 3.015  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__mux4_1
