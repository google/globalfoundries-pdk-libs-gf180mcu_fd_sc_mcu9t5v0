* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__xor3_4 A1 A2 A3 Z VDD VNW VPW VSS
*.PININFO A1:I A2:I A3:I Z:O VDD:P VNW:P VPW:P VSS:G
*.EQN Z=!((!((A1 * A2) + !(A1 + A2)) * A3) + !(!((A1 * A2) + !(A1 + A2)) + A3))
M_i_14 I A2 VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_15 VSS A1 I VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_2 I2 I VSS VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_0 net_0 A1 I2 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_1 VSS A2 net_0 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_18 net_5 I2 I3 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_19 VSS A3 net_5 VPW nmos_5p0 W=0.360000U L=0.600000U
M_i_10 net_2 I3 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_8 Z_neg A3 net_2 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_9 net_2 I2 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_3 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_2 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_1 VSS Z_neg Z VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_6_0 Z Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_16 net_4 A2 I VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_17 VDD A1 net_4 VNW pmos_5p0 W=0.360000U L=0.500000U
M_i_5 net_1 I VDD VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_3 I2 A1 net_1 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_4 net_1 A2 I2 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_20 I3 I2 VDD VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_21 VDD A3 I3 VNW pmos_5p0 W=0.495000U L=0.500000U
M_i_13 Z_neg I3 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_11 net_3 A3 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_12 VDD I2 net_3 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_3 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_2 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_1 VDD Z_neg Z VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_7_0 Z Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
