# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.353 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2 0.97 2 0.97 3.27 0.63 3.27  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.5506 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.665 3.96 2.88 3.96 2.88 1.215 2.33 1.215 2.33 0.71 3.11 0.71 3.11 4.3 2.665 4.3  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.96 1.495 3.96 1.495 4.59 2.65 4.59 3.685 4.59 3.685 3.55 3.915 3.55 3.915 4.59 4.48 4.59 4.48 5.49 2.65 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 4.015 0.45 4.015 1.215 3.785 1.215 3.785 0.45 1.595 0.45 1.595 1.215 1.365 1.215 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 3.5 1.37 3.5 1.37 1.77 0.245 1.77 0.245 0.875 0.475 0.875 0.475 1.54 1.6 1.54 1.6 2.27 2.65 2.27 2.65 2.5 1.6 2.5 1.6 3.73 0.475 3.73 0.475 4.36 0.245 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_2
