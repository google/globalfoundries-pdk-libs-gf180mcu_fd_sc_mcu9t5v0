# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__icgtn_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__icgtn_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.16 BY 5.04 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.64 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.35 1.77 11.61 1.77 11.61 2.71 11.35 2.71  ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.345 1.82 2.65 1.82 2.65 3.27 2.345 3.27  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.11 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 1.77 0.97 1.77 0.97 2.71 0.71 2.71  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.9432 ;
    PORT
      LAYER METAL1 ;
        POLYGON 16.03 2.69 17.51 2.69 18.07 2.69 18.07 1.6 16.03 1.6 16.03 0.79 16.31 0.79 16.31 1.3 18.32 1.3 18.32 0.79 18.55 0.79 18.55 3.96 18.07 3.96 18.07 2.92 17.51 2.92 16.26 2.92 16.26 3.96 16.03 3.96  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.325 4.59 1.325 3.15 1.555 3.15 1.555 4.59 2.715 4.59 5.82 4.59 5.82 3.15 6.05 3.15 6.05 4.59 8.25 4.59 8.58 4.59 8.58 3.15 8.81 3.15 8.81 4.59 9.305 4.59 12.08 4.59 12.08 3.785 12.31 3.785 12.31 4.59 12.75 4.59 15.01 4.59 15.01 3.15 15.24 3.15 15.24 4.59 17.05 4.59 17.05 3.15 17.28 3.15 17.28 4.59 17.51 4.59 19.09 4.59 19.09 3.15 19.32 3.15 19.32 4.59 20.16 4.59 20.16 5.49 17.51 5.49 12.75 5.49 9.305 5.49 8.25 5.49 2.715 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 20.16 -0.45 20.16 0.45 19.67 0.45 19.67 1.6 19.44 1.6 19.44 0.45 17.43 0.45 17.43 1.07 17.2 1.07 17.2 0.45 15.19 0.45 15.19 1.6 14.96 1.6 14.96 0.45 14.45 0.45 14.45 1.13 14.22 1.13 14.22 0.45 12.21 0.45 12.21 1.13 11.98 1.13 11.98 0.45 8.81 0.45 8.81 1.13 8.58 1.13 8.58 0.45 5.81 0.45 5.81 1.13 5.58 1.13 5.58 0.45 1.65 0.45 1.65 1.075 1.31 1.075 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.79 0.475 0.79 0.475 1.305 2.485 1.305 2.485 0.79 2.715 0.79 2.715 1.535 0.245 1.535  ;
        POLYGON 3.405 1.845 6.7 1.845 6.7 0.79 7.07 0.79 7.07 3.9 6.84 3.9 6.84 2.075 4.81 2.075 4.81 2.46 4.47 2.46 4.47 2.075 3.405 2.075  ;
        POLYGON 3.175 2.565 4.265 2.565 4.265 2.69 6.51 2.69 6.51 4.13 8.02 4.13 8.02 1.82 8.25 1.82 8.25 4.36 6.28 4.36 6.28 2.92 4.29 2.92 4.29 3.96 4.06 3.96 4.06 2.795 2.945 2.795 2.945 1.385 3.62 1.385 3.62 0.79 3.85 0.79 3.85 1.615 3.175 1.615  ;
        POLYGON 7.46 0.79 7.69 0.79 7.69 1.36 8.71 1.36 8.71 1.875 9.305 1.875 9.305 2.105 8.48 2.105 8.48 1.59 7.79 1.59 7.79 3.9 7.46 3.9  ;
        POLYGON 10.36 1.23 11.09 1.23 11.09 2.935 11.29 2.935 11.29 3.275 10.86 3.275 10.86 1.46 10.59 1.46 10.59 2.2 10.36 2.2  ;
        POLYGON 9.6 0.79 9.93 0.79 9.93 3.505 11.63 3.505 11.63 3.325 12.52 3.325 12.52 2.475 12.75 2.475 12.75 3.555 11.855 3.555 11.855 3.735 9.83 3.735 9.83 3.96 9.6 3.96  ;
        POLYGON 13.045 1.285 13.385 1.285 13.385 1.305 14.07 1.305 14.07 1.98 17.51 1.98 17.51 2.32 14.07 2.32 14.07 3.96 13.84 3.96 13.84 1.535 13.045 1.535  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__icgtn_4
