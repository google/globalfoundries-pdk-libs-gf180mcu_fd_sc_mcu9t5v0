# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi222_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 26.32 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.865 1.755 25.095 1.755 25.095 2.555 24.865 2.555 24.865 1.985 21.015 1.985 21.015 2.4 20.785 2.4 20.785 1.985 19.45 1.985 19.45 2.15 18.095 2.15 18.095 2.555 17.865 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.75 2.27 20.32 2.27 20.32 2.63 22.595 2.63 22.595 2.215 23.055 2.215 23.055 2.77 22.78 2.77 22.78 2.86 20.135 2.86 20.135 2.77 19.75 2.77  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.67 1.37 12.775 1.37 12.775 1.425 16.835 1.425 16.835 2.555 16.605 2.555 16.605 1.655 12.855 1.655 12.855 2.4 12.625 2.4 12.625 1.6 9.93 1.6 9.93 2.555 9.67 2.555  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.69 1.83 12.33 1.83 12.33 2.63 13.955 2.63 13.955 2.54 14.665 2.54 14.665 2.215 14.895 2.215 14.895 2.77 14.14 2.77 14.14 2.86 12.1 2.86 12.1 2.5 11.69 2.5  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.755 8.055 1.755 8.055 2.555 7.825 2.555 7.825 2.15 6.31 2.15 6.31 1.985 3.975 1.985 3.975 2.555 3.745 2.555 3.745 1.985 1.055 1.985 1.055 2.555 0.825 2.555  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.215 3.515 2.215 3.515 2.785 5.49 2.785 5.49 2.625 5.785 2.625 5.785 2.215 6.015 2.215 6.015 2.855 5.71 2.855 5.71 3.015 3.285 3.015 3.285 2.445 2.09 2.445 2.09 2.71 1.83 2.71  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.2844 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.19 0.91 13.49 0.91 13.49 0.925 24.73 0.925 24.73 0.71 25.73 0.71 25.73 1.195 17.515 1.195 17.515 2.785 17.895 2.785 17.895 3 19.925 3 19.925 3.09 23.035 3.09 23.035 3 24.655 3 24.655 3.9 24.425 3.9 24.425 3.23 23.22 3.23 23.22 3.32 22.615 3.32 22.615 3.9 22.385 3.9 22.385 3.32 20.575 3.32 20.575 3.9 20.345 3.9 20.345 3.32 19.74 3.32 19.74 3.23 18.535 3.23 18.535 3.9 18.305 3.9 18.305 3.23 17.665 3.23 17.665 3.015 17.285 3.015 17.285 1.155 13.405 1.155 13.405 1.14 8.69 1.14 8.69 1.195 0.19 1.195  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.245 0.475 3.245 0.475 4.59 2.285 4.59 2.285 3.705 2.515 3.705 2.515 4.59 4.325 4.59 4.325 3.705 4.555 3.705 4.555 4.59 6.365 4.59 6.365 3.56 6.595 3.56 6.595 4.59 8.405 4.59 8.405 3.545 8.635 3.545 8.635 4.59 25.675 4.59 26.32 4.59 26.32 5.49 25.675 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 26.32 -0.45 26.32 0.45 23.635 0.45 23.635 0.695 23.405 0.695 23.405 0.45 19.555 0.45 19.555 0.695 19.325 0.695 19.325 0.45 15.475 0.45 15.475 0.695 15.245 0.695 15.245 0.45 11.45 0.45 11.45 0.68 11.11 0.68 11.11 0.45 6.65 0.45 6.65 0.68 6.31 0.68 6.31 0.45 2.57 0.45 2.57 0.68 2.23 0.68 2.23 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 3.245 5.93 3.245 5.93 3.085 9.455 3.085 9.455 3.09 14.325 3.09 14.325 3 16.495 3 16.495 3.9 16.265 3.9 16.265 3.23 14.51 3.23 14.51 3.9 14.225 3.9 14.225 3.32 12.415 3.32 12.415 3.9 12.185 3.9 12.185 3.32 10.375 3.32 10.375 3.9 10.145 3.9 10.145 3.32 9.405 3.32 9.405 3.315 7.615 3.315 7.615 4.055 7.385 4.055 7.385 3.315 6.15 3.315 6.15 3.475 5.575 3.475 5.575 4.055 5.345 4.055 5.345 3.475 3.535 3.475 3.535 4.055 3.305 4.055 3.305 3.475 1.495 3.475 1.495 4.055 1.265 4.055  ;
        POLYGON 9.125 3.545 9.355 3.545 9.355 4.13 11.165 4.13 11.165 3.55 11.395 3.55 11.395 4.13 13.205 4.13 13.205 3.55 13.435 3.55 13.435 4.13 15.245 4.13 15.245 3.46 15.475 3.46 15.475 4.13 17.285 4.13 17.285 3.405 17.515 3.405 17.515 4.13 19.325 4.13 19.325 3.46 19.555 3.46 19.555 4.13 21.365 4.13 21.365 3.55 21.595 3.55 21.595 4.13 23.405 4.13 23.405 3.46 23.635 3.46 23.635 4.13 25.445 4.13 25.445 3.245 25.675 3.245 25.675 4.36 9.125 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi222_4
