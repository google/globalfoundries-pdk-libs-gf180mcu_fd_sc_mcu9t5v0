# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dlya_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlya_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.16 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.77 1.045 1.77 1.045 2.495 0.705 2.495  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 4.07 5.185 4.07 5.535 4.07 5.535 0.845 5.865 0.845 5.865 4.33 5.185 4.33 5.13 4.33  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.24 1.495 3.24 1.495 4.59 2.035 4.59 4.125 4.59 4.125 3.24 4.355 3.24 4.355 4.59 5.185 4.59 6.16 4.59 6.16 5.49 5.185 5.49 2.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.16 -0.45 6.16 0.45 4.745 0.45 4.745 0.695 4.515 0.695 4.515 0.45 1.595 0.45 1.595 1.62 1.365 1.62 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.28 0.475 1.28 0.475 2.725 1.805 2.725 1.805 1.74 2.035 1.74 2.035 2.955 0.475 2.955 0.475 3.58 0.245 3.58  ;
        POLYGON 2.385 1.28 2.715 1.28 2.715 1.795 3.83 1.795 3.83 2.495 2.615 2.495 2.615 3.58 2.385 3.58  ;
        POLYGON 3.105 2.78 4.06 2.78 4.06 1.745 4.055 1.745 4.055 0.91 3 0.91 3 0.68 4.285 0.68 4.285 1.695 5.185 1.695 5.185 2.585 4.29 2.585 4.29 3.01 3.335 3.01 3.335 3.58 3.105 3.58  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlya_1
