# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai211_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.6 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 2.27 2.17 2.27 2.17 2.71 1.83 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.215 1.015 2.215 1.015 2.71 0.71 2.71  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 2.27 3.29 2.27 3.29 2.71 2.95 2.71  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.522 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.99 2.27 4.33 2.27 4.33 2.71 3.99 2.71  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.4988 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 1.14 1.595 1.14 1.595 3.09 2.715 3.09 4.835 3.09 4.835 4.36 4.605 4.36 4.605 3.32 2.715 3.32 2.615 3.32 2.615 4.36 2.385 4.36 2.385 3.32 1.27 3.32  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 3.55 0.575 3.55 0.575 4.59 2.715 4.59 3.585 4.59 3.585 3.55 3.815 3.55 3.815 4.59 5.6 4.59 5.6 5.49 2.715 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 5.6 -0.45 5.6 0.45 4.835 0.45 4.835 1.655 4.605 1.655 4.605 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.68 2.715 0.68 2.715 1.655 2.485 1.655 2.485 0.91 0.475 0.91 0.475 1.655 0.245 1.655  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai211_1
