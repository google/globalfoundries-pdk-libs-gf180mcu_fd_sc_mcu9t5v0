# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.92 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.5 1.77 3.77 1.77 3.77 2.72 3.5 2.72  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 1.31 4.26 1.31 4.26 1.355 5.19 1.355 5.19 1.21 5.45 1.21 5.45 1.92 5.87 1.92 5.87 2.72 5.64 2.72 5.64 2.15 5.19 2.15 5.19 1.585 4.35 1.585 4.35 2.72 4.12 2.72 4.12 1.54 0.97 1.54 0.97 2.72 0.74 2.72  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.34 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 1.77 2.65 1.77 2.65 2.72 2.39 2.72  ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.035 0.785 14.41 0.785 14.41 1.825 16.325 1.825 16.325 0.785 16.555 0.785 16.555 2.055 14.41 2.055 14.41 3.415 16.305 3.415 16.305 4.36 16.075 4.36 16.075 3.645 14.265 3.645 14.265 4.36 14.035 4.36  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.32 4.59 1.32 3.55 1.55 3.55 1.55 4.59 3.24 4.59 3.24 3.87 3.47 3.87 3.47 4.59 7.61 4.59 7.61 3.7 7.84 3.7 7.84 4.59 9.88 4.59 9.88 3.55 10.11 3.55 10.11 4.59 10.84 4.59 12.07 4.59 12.07 3.55 12.3 3.55 12.3 4.59 13.015 4.59 13.015 3.875 13.245 3.875 13.245 4.59 13.74 4.59 15.055 4.59 15.055 3.875 15.285 3.875 15.285 4.59 17.095 4.59 17.095 3.875 17.325 3.875 17.325 4.59 17.92 4.59 17.92 5.49 13.74 5.49 10.84 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 17.92 -0.45 17.92 0.45 17.675 0.45 17.675 1.595 17.445 1.595 17.445 0.45 15.435 0.45 15.435 1.595 15.205 1.595 15.205 0.45 13.195 0.45 13.195 1.595 12.965 1.595 12.965 0.45 12.45 0.45 12.45 1.125 12.22 1.125 12.22 0.45 10.21 0.45 10.21 1.125 9.98 1.125 9.98 0.45 7.97 0.45 7.97 1.125 7.74 1.125 7.74 0.45 1.685 0.45 1.685 1.07 1.345 1.07 1.345 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.28 0.785 0.51 0.785 0.51 2.95 5.04 2.95 5.04 2.38 5.27 2.38 5.27 3.18 0.53 3.18 0.53 4.36 0.28 4.36  ;
        POLYGON 2.22 3.41 5.55 3.41 5.55 3.81 6.1 3.81 6.1 0.98 4.81 0.98 4.81 1.125 4.58 1.125 4.58 0.75 6.33 0.75 6.33 1.92 8.46 1.92 8.46 2.72 8.23 2.72 8.23 2.15 6.33 2.15 6.33 4.04 5.32 4.04 5.32 3.64 2.45 3.64 2.45 4.04 2.22 4.04  ;
        POLYGON 7.17 2.38 7.4 2.38 7.4 2.95 8.86 2.95 8.86 0.785 9.09 0.785 9.09 2.95 10.61 2.95 10.61 2.38 10.84 2.38 10.84 3.18 9.04 3.18 9.04 4.36 8.81 4.36 8.81 3.18 7.17 3.18  ;
        POLYGON 11.05 3.55 11.095 3.55 11.095 0.785 11.33 0.785 11.33 2.435 13.74 2.435 13.74 2.665 11.325 2.665 11.325 4.36 11.05 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_4
