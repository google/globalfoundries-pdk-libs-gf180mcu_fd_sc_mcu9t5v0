# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai221_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 24.08 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 15.03 2.27 15.37 2.27 15.37 3.04 19.14 3.04 19.14 2.215 19.37 2.215 19.37 2.89 20.96 2.89 20.96 2.27 22.97 2.27 22.97 2.5 21.19 2.5 21.19 3.27 15.03 3.27  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 17.27 2.27 17.51 2.27 17.51 1.755 19.83 1.755 19.83 2.27 20.73 2.27 20.73 2.5 19.6 2.5 19.6 1.985 17.77 1.985 17.77 2.5 17.27 2.5  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.87 2.27 1.21 2.27 1.21 2.73 4.07 2.73 4.07 2.27 4.41 2.27 4.41 2.73 6.85 2.73 6.85 2.27 8.86 2.27 8.86 2.5 7.08 2.5 7.08 2.96 0.87 2.96  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.828 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.06 2.27 3.4 2.27 3.4 2.02 3.46 2.02 3.46 1.77 4.87 1.77 4.87 2.27 6.62 2.27 6.62 2.5 4.64 2.5 4.64 2.04 3.86 2.04 3.86 2.175 3.63 2.175 3.63 2.5 3.06 2.5  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.088 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.99 2.27 13.515 2.27 13.57 2.27 13.57 2.71 13.515 2.71 10.99 2.71  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.615 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.345 3.19 4.905 3.19 4.905 3.5 13.515 3.5 23.2 3.5 23.2 1.97 20.06 1.97 20.06 1.52 15.525 1.52 15.525 1.14 15.755 1.14 15.755 1.29 17.71 1.29 17.71 1.14 18.05 1.14 18.05 1.29 20.005 1.29 20.005 1.14 20.29 1.14 20.29 1.74 22.245 1.74 22.245 1.14 22.475 1.14 22.475 1.74 23.495 1.74 23.495 4.36 23.265 4.36 23.265 3.73 19.065 3.73 19.065 4.36 18.57 4.36 18.57 3.73 14.535 3.73 14.535 4.36 14.305 4.36 14.305 3.73 13.515 3.73 12.395 3.73 12.395 4.36 12.165 4.36 12.165 3.73 9.385 3.73 9.385 4.36 9.155 4.36 9.155 3.73 4.905 3.73 4.905 4.36 4.675 4.36 4.675 3.42 0.575 3.42 0.575 4.36 0.345 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.65 2.665 3.65 2.665 4.59 6.915 4.59 6.915 3.96 7.145 3.96 7.145 4.59 10.945 4.59 10.945 3.96 11.175 3.96 11.175 4.59 13.185 4.59 13.185 3.96 13.415 3.96 13.415 4.59 13.515 4.59 16.595 4.59 16.595 3.96 16.825 3.96 16.825 4.59 21.075 4.59 21.075 3.96 21.305 3.96 21.305 4.59 23.595 4.59 24.08 4.59 24.08 5.49 23.595 5.49 13.515 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 24.08 -0.45 24.08 0.45 9.435 0.45 9.435 1.04 9.205 1.04 9.205 0.45 7.195 0.45 7.195 1.04 6.965 1.04 6.965 0.45 4.955 0.45 4.955 1.04 4.725 1.04 4.725 0.45 2.715 0.45 2.715 1.51 2.485 1.51 2.485 0.45 0.475 0.45 0.475 1.51 0.245 1.51 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.365 0.7 1.595 0.7 1.595 1.74 2.945 1.74 2.945 1.28 3.605 1.28 3.605 0.7 3.835 0.7 3.835 1.28 5.845 1.28 5.845 0.7 6.075 0.7 6.075 1.28 8.085 1.28 8.085 0.7 8.315 0.7 8.315 1.28 10.99 1.28 10.99 1.14 11.33 1.14 11.33 1.28 13.285 1.28 13.285 1.14 13.515 1.14 13.515 1.51 3.175 1.51 3.175 1.97 1.365 1.97  ;
        POLYGON 9.925 0.68 23.595 0.68 23.595 1.51 23.365 1.51 23.365 0.91 21.355 0.91 21.355 1.51 21.125 1.51 21.125 0.91 19.17 0.91 19.17 0.985 18.83 0.985 18.83 0.91 16.93 0.91 16.93 0.985 16.59 0.985 16.59 0.91 14.69 0.91 14.69 0.985 14.35 0.985 14.35 0.91 12.45 0.91 12.45 0.985 12.11 0.985 12.11 0.91 10.155 0.91 10.155 1.04 9.925 1.04  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai221_4
