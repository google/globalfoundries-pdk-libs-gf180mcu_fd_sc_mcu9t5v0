# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__clkbuf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 28 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.824 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 2.125 7.965 2.125 7.965 2.84 0.685 2.84  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 12.4048 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.505 3.09 17.105 3.09 17.985 3.09 17.985 1.895 10.505 1.895 10.505 0.945 10.735 0.945 10.735 1.515 12.745 1.515 12.745 0.945 12.975 0.945 12.975 1.665 14.985 1.665 14.985 0.945 15.215 0.945 15.215 1.665 17.225 1.665 17.225 0.945 17.455 0.945 17.455 1.515 19.465 1.515 19.465 0.945 19.695 0.945 19.695 1.515 21.705 1.515 21.705 0.945 21.935 0.945 21.935 1.515 23.945 1.515 23.945 0.945 24.175 0.945 24.175 1.515 26.185 1.515 26.185 0.945 26.415 0.945 26.415 1.745 18.735 1.745 18.735 3.09 26.245 3.09 26.315 3.09 26.315 4.36 26.245 4.36 26.085 4.36 26.085 3.32 24.075 3.32 24.075 4.36 23.845 4.36 23.845 3.32 21.835 3.32 21.835 4.36 21.605 4.36 21.605 3.32 19.595 3.32 19.595 4.36 19.365 4.36 19.365 3.32 17.355 3.32 17.355 4.36 17.125 4.36 17.125 3.32 17.105 3.32 15.115 3.32 15.115 4.36 14.885 4.36 14.885 3.32 12.875 3.32 12.875 4.36 12.645 4.36 12.645 3.32 10.735 3.32 10.735 4.36 10.505 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 9.105 4.59 9.105 3.875 9.335 3.875 9.335 4.59 11.525 4.59 11.525 3.55 11.755 3.55 11.755 4.59 13.765 4.59 13.765 3.55 13.995 3.55 13.995 4.59 16.005 4.59 16.005 3.55 16.235 3.55 16.235 4.59 17.105 4.59 18.245 4.59 18.245 3.55 18.475 3.55 18.475 4.59 20.485 4.59 20.485 3.55 20.715 3.55 20.715 4.59 22.725 4.59 22.725 3.55 22.955 3.55 22.955 4.59 24.965 4.59 24.965 3.55 25.195 3.55 25.195 4.59 26.245 4.59 27.205 4.59 27.205 3.55 27.435 3.55 27.435 4.59 28 4.59 28 5.49 26.245 5.49 17.105 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 28 -0.45 28 0.45 27.535 0.45 27.535 1.285 27.305 1.285 27.305 0.45 25.295 0.45 25.295 1.215 25.065 1.215 25.065 0.45 23.055 0.45 23.055 1.215 22.825 1.215 22.825 0.45 20.815 0.45 20.815 1.285 20.585 1.285 20.585 0.45 18.575 0.45 18.575 1.215 18.345 1.215 18.345 0.45 16.335 0.45 16.335 1.215 16.105 1.215 16.105 0.45 14.095 0.45 14.095 1.285 13.865 1.285 13.865 0.45 11.855 0.45 11.855 1.285 11.625 1.285 11.625 0.45 9.435 0.45 9.435 1.285 9.205 1.285 9.205 0.45 7.195 0.45 7.195 1.285 6.965 1.285 6.965 0.45 4.955 0.45 4.955 1.285 4.725 1.285 4.725 0.45 2.715 0.45 2.715 1.285 2.485 1.285 2.485 0.45 0.475 0.45 0.475 1.285 0.245 1.285 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 3.09 8.32 3.09 8.32 1.745 1.365 1.745 1.365 0.945 1.595 0.945 1.595 1.515 3.605 1.515 3.605 0.945 3.835 0.945 3.835 1.515 5.845 1.515 5.845 0.945 6.075 0.945 6.075 1.515 8.085 1.515 8.085 0.945 8.55 0.945 8.55 2.215 17.105 2.215 17.105 2.555 8.55 2.555 8.55 4.36 8.085 4.36 8.085 3.32 5.975 3.32 5.975 4.36 5.745 4.36 5.745 3.32 3.735 3.32 3.735 4.36 3.505 4.36 3.505 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
        POLYGON 18.965 2.215 26.245 2.215 26.245 2.555 18.965 2.555  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__clkbuf_16
