# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai222_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 15.12 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 10.605 2.215 10.835 2.215 10.835 2.94 12.27 2.94 12.27 2.215 14.005 2.215 14.005 2.71 12.5 2.71 12.5 3.17 10.605 3.17  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.35 2.215 11.715 2.215 11.715 2.71 11.35 2.71  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.19 2.215 6.165 2.215 6.165 3.04 9.035 3.04 9.295 3.04 9.295 2.215 9.525 2.215 9.525 3.27 9.035 3.27 5.19 3.27  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.87 2.215 7.285 2.215 7.285 2.71 6.87 2.71  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.925 2.215 1.155 2.215 1.155 2.785 4.07 2.785 4.07 1.77 4.33 1.77 4.33 3.015 0.925 3.015  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.555 1.83 2.555  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.57 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.345 3.32 4.9 3.32 4.9 3.5 8.87 3.5 8.87 4.13 9.035 4.13 9.875 4.13 9.875 3.4 14.355 3.4 14.355 1.95 11.045 1.95 11.045 1.14 11.275 1.14 11.275 1.72 13.285 1.72 13.285 1.14 13.515 1.14 13.515 1.72 14.585 1.72 14.585 4.36 14.355 4.36 14.355 3.63 10.105 3.63 10.105 4.36 9.035 4.36 8.49 4.36 8.49 3.73 4.905 3.73 4.905 4.36 4.675 4.36 4.675 3.55 0.575 3.55 0.575 4.36 0.345 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.78 2.665 3.78 2.665 4.59 7.635 4.59 7.635 3.96 7.865 3.96 7.865 4.59 9.035 4.59 12.115 4.59 12.115 3.86 12.345 3.86 12.345 4.59 14.635 4.59 15.12 4.59 15.12 5.49 14.635 5.49 9.035 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 15.12 -0.45 15.12 0.45 4.955 0.45 4.955 0.695 4.725 0.695 4.725 0.45 2.715 0.45 2.715 0.695 2.485 0.695 2.485 0.45 0.475 0.45 0.475 1.655 0.245 1.655 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.365 0.73 1.595 0.73 1.595 0.925 3.605 0.925 3.605 0.73 3.835 0.73 3.835 1.14 9.035 1.14 9.035 1.54 1.365 1.54  ;
        POLYGON 5.39 0.68 14.635 0.68 14.635 1.49 14.405 1.49 14.405 0.91 12.395 0.91 12.395 1.49 12.165 1.49 12.165 0.91 10.155 0.91 10.155 1.575 9.925 1.575 9.925 0.91 5.39 0.91  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai222_2
