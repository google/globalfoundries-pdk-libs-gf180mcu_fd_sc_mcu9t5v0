# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__tiel
  CLASS core gf180mcu_fd_sc_mcu9t5v0__tielOW ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__tiel 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 2.24 BY 5.04 ;
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.2904 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.215 1.21 1.595 1.21 1.595 1.59 1.215 1.59  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.345 4.59 0.345 2.945 0.575 2.945 0.575 4.59 1.595 4.59 2.24 4.59 2.24 5.49 1.595 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 2.24 -0.45 2.24 0.45 0.475 0.45 0.475 1.355 0.245 1.355 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.87 2.47 1.595 2.47 1.595 3.685 1.365 3.685 1.365 2.7 0.87 2.7  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__tiel
