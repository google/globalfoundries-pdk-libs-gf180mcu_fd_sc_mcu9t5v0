# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__oai21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__oai21_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 4.48 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.77 2.09 1.77 2.09 2.555 1.83 2.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.68 2.27 1.02 2.27 1.02 2.71 0.68 2.71  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.6145 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.95 2.27 3.29 2.27 3.29 2.71 2.95 2.71  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9119 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.27 1.14 1.595 1.14 1.595 2.785 2.615 2.785 2.615 4.36 2.385 4.36 2.385 3.015 1.27 3.015  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.295 4.59 0.295 3.55 0.525 3.55 0.525 4.59 2.715 4.59 3.585 4.59 3.585 3.55 3.815 3.55 3.815 4.59 4.48 4.59 4.48 5.49 2.715 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 4.48 -0.45 4.48 0.45 3.835 0.45 3.835 1.655 3.605 1.655 3.605 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.68 2.715 0.68 2.715 1.655 2.485 1.655 2.485 0.91 0.475 0.91 0.475 1.655 0.245 1.655  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__oai21_1
