# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__addh_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__addh_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.285 2.215 2.515 2.215 2.515 2.95 5.845 2.95 5.845 2.215 6.075 2.215 6.075 3.27 2.285 3.27  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.707 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.95 2.27 5.195 2.27 5.195 2.65 2.95 2.65  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 0.845 0.575 0.845 0.575 4.36 0.15 4.36  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 8.55 1.21 8.945 1.21 8.945 0.845 9.175 0.845 9.175 4.36 8.845 4.36 8.845 1.59 8.55 1.59  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.55 1.595 3.55 1.595 4.59 3.645 4.59 3.645 3.96 3.875 3.96 3.875 4.59 4.385 4.59 4.385 3.96 4.615 3.96 4.615 4.59 7.645 4.59 7.645 3.55 7.875 3.55 7.875 4.59 8.495 4.59 9.52 4.59 9.52 5.49 8.495 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 7.875 0.45 7.875 1.355 7.645 1.355 7.645 0.45 1.595 0.45 1.595 1.35 1.365 1.35 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 4.285 0.68 6.755 0.68 6.755 1.355 6.525 1.355 6.525 0.91 4.515 0.91 4.515 1.355 4.285 1.355  ;
        POLYGON 2.055 3.5 6.725 3.5 6.725 2.27 7.35 2.27 7.35 2.5 6.955 2.5 6.955 3.73 2.855 3.73 2.855 4.36 2.625 4.36 2.625 3.73 1.825 3.73 1.825 2.555 0.925 2.555 0.925 2.215 1.825 2.215 1.825 1.07 3.85 1.07 3.85 1.3 2.055 1.3  ;
        POLYGON 6.57 3.96 7.185 3.96 7.185 3.09 7.58 3.09 7.58 1.985 5.405 1.985 5.405 1.14 5.635 1.14 5.635 1.755 7.81 1.755 7.81 2.215 8.495 2.215 8.495 2.555 7.81 2.555 7.81 3.32 7.415 3.32 7.415 4.19 6.57 4.19  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__addh_1
