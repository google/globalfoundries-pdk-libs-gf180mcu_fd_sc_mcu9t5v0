# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dlya_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dlya_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.035 1.05 2.035 1.05 2.735 0.71 2.735  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.68 2.95 7.115 2.95 7.345 2.95 7.345 2.04 5.63 2.04 5.63 0.77 5.86 0.77 5.86 1.81 7.87 1.81 7.87 0.77 8.1 0.77 8.1 2.04 7.575 2.04 7.575 2.98 8.05 2.98 8.05 4.25 7.82 4.25 7.82 3.21 7.115 3.21 5.91 3.21 5.91 4.25 5.68 4.25  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.27 4.59 1.27 3.44 1.5 3.44 1.5 4.59 2.095 4.59 4.28 4.59 4.28 3.44 4.51 3.44 4.51 4.59 6.7 4.59 6.7 3.44 6.93 3.44 6.93 4.59 7.115 4.59 8.89 4.59 8.89 3.44 9.12 3.44 9.12 4.59 9.52 4.59 9.52 5.49 7.115 5.49 2.095 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 9.22 0.45 9.22 1.58 8.99 1.58 8.99 0.45 6.98 0.45 6.98 1.58 6.75 1.58 6.75 0.45 4.56 0.45 4.56 1.11 4.33 1.11 4.33 0.45 1.6 0.45 1.6 1.11 1.37 1.11 1.37 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.25 0.77 0.48 0.77 0.48 2.965 1.755 2.965 1.755 2.035 2.095 2.035 2.095 3.195 0.48 3.195 0.48 3.78 0.25 3.78  ;
        POLYGON 2.39 2.505 3.7 2.505 3.7 2.03 2.49 2.03 2.49 0.77 2.72 0.77 2.72 1.8 3.985 1.8 3.985 2.735 2.62 2.735 2.62 3.78 2.39 3.78  ;
        POLYGON 3.26 2.98 4.215 2.98 4.215 1.57 3.21 1.57 3.21 0.77 3.44 0.77 3.44 1.34 4.445 1.34 4.445 2.27 7.115 2.27 7.115 2.5 4.445 2.5 4.445 3.21 3.49 3.21 3.49 3.78 3.26 3.78  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dlya_4
