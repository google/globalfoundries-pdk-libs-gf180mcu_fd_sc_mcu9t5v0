* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__tieh Z VDD VNW VPW VSS
*.PININFO Z:O VDD:P VNW:P VPW:P VSS:G
M_n_tran_1 VSS A A VPW nmos_5p0 W=0.660000U L=0.600000U
M_p_tran_2 VDD A Z VNW pmos_5p0 W=0.900000U L=0.500000U
.ENDS
