* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4 D RN CLKN Q VDD VNW VPW VSS
*.PININFO D:I RN:I CLKN:I Q:O VDD:P VNW:P VPW:P VSS:G
M_tn13 ncki CLKN VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn10 cki ncki VSS VPW nmos_5p0 W=0.790000U L=0.600000U
M_tn11 net6 D VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn15 net6 cki net1 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn14 net1 ncki net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn8 net12 net2 net15 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn9 VSS RN net12 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn18 VSS net1 net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn0 net8 ncki net2 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn1 net11 cki net8 VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn12 net11 net4 VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn5 net0 RN VSS VPW nmos_5p0 W=0.700000U L=0.600000U
M_tn4 net4 net8 net0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_42 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_42_63 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tn3_69 Q net4 VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_tp11 ncki CLKN VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp8 cki ncki VDD VNW pmos_5p0 W=1.380000U L=0.500000U
M_tp9 VDD D net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp15 net1 ncki net6 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp7 net9 cki net1 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp6 VDD net2 net9 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp12 net9 RN VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp18 VDD net1 net2 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp2 net2 cki net8 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp3 net8 ncki net11 VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp10 net11 net4 VDD VNW pmos_5p0 W=1.000000U L=0.500000U
M_tp5 net4 RN VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp4 VDD net8 net4 VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_40 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_40_64 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_tp1_66 Q net4 VDD VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
