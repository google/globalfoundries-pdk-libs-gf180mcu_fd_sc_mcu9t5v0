# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__latrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__latrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 12.88 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER METAL1 ;
        POLYGON 2.95 1.77 3.295 1.77 3.295 2.71 2.95 2.71  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 2.084 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.705 1.21 0.97 1.21 0.97 1.31 3.905 1.31 3.905 1.495 5.195 1.495 5.195 2.44 5.5 2.44 5.5 2.67 4.965 2.67 4.965 1.725 4.135 1.725 4.135 2.295 3.675 2.295 3.675 1.54 0.97 1.54 0.97 2.295 0.705 2.295  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.34 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.83 1.77 2.455 1.77 2.455 2.71 1.83 2.71  ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.386 ;
    PORT
      LAYER METAL1 ;
        POLYGON 11.91 0.845 12.355 0.845 12.355 4.36 11.91 4.36  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.265 4.59 1.265 3.55 1.495 3.55 1.495 4.59 3.025 4.59 3.025 3.86 3.255 3.86 3.255 4.59 6.63 4.59 6.63 3.55 6.86 3.55 6.86 4.59 9.215 4.59 9.215 3.55 9.445 3.55 9.445 4.59 9.835 4.59 11.055 4.59 11.055 3.875 11.285 3.875 11.285 4.59 11.62 4.59 12.88 4.59 12.88 5.49 11.62 5.49 9.835 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 12.88 -0.45 12.88 0.45 11.235 0.45 11.235 1.605 11.005 1.605 11.005 0.45 9.395 0.45 9.395 1.135 9.165 1.135 9.165 0.45 7.375 0.45 7.375 1.135 7.145 1.135 7.145 0.45 1.65 0.45 1.65 1.08 1.31 1.08 1.31 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 0.795 0.475 0.795 0.475 2.94 4.505 2.94 4.505 1.955 4.735 1.955 4.735 3.17 0.475 3.17 0.475 4.36 0.245 4.36  ;
        POLYGON 2.005 3.4 5.015 3.4 5.015 4.13 5.73 4.13 5.73 1.495 6.45 1.495 6.45 1.135 4.345 1.135 4.345 0.795 6.68 0.795 6.68 1.535 7.78 1.535 7.78 2.295 7.55 2.295 7.55 1.765 6.55 1.765 6.55 1.725 5.96 1.725 5.96 4.36 4.785 4.36 4.785 3.63 2.235 3.63 2.235 4.36 2.005 4.36  ;
        POLYGON 6.19 1.955 6.42 1.955 6.42 2.525 8.01 2.525 8.01 2.065 8.445 2.065 8.445 0.795 8.675 0.795 8.675 1.955 9.835 1.955 9.835 2.295 8.24 2.295 8.24 4.36 7.83 4.36 7.83 2.755 6.19 2.755  ;
        POLYGON 10.235 1.225 10.515 1.225 10.515 2.03 11.62 2.03 11.62 2.26 10.465 2.26 10.465 4.36 10.235 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__latrnq_1
