# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__aoi211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__aoi211_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 9.52 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.765 1.77 2.955 1.77 2.955 2.215 1.765 2.215  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.252 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.63 2.305 1.155 2.305 1.155 2.445 3.51 2.445 3.51 1.77 3.77 1.77 3.77 2.775 0.63 2.775  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER METAL1 ;
        POLYGON 4.56 1.725 5.45 1.725 5.45 2.47 8.43 2.47 8.43 2.7 4.56 2.7  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.778 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.75 1.77 7.295 1.77 7.295 2.15 5.75 2.15  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.341 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.21 3.4 4.07 3.4 4.07 1.525 2.205 1.525 2.205 0.715 2.435 0.715 2.435 1.265 4.73 1.265 4.73 0.93 5.465 0.93 5.465 0.695 5.695 0.695 5.695 0.93 7.705 0.93 7.705 0.79 7.935 0.79 7.935 1.16 4.96 1.16 4.96 1.495 4.33 1.495 4.33 3.63 1.21 3.63  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 6.505 4.59 6.505 4.345 6.735 4.345 6.735 4.59 8.815 4.59 9.52 4.59 9.52 5.49 8.815 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 9.52 -0.45 9.52 0.45 9.055 0.45 9.055 0.7 8.825 0.7 8.825 0.45 6.815 0.45 6.815 0.7 6.585 0.7 6.585 0.45 4.395 0.45 4.395 0.7 4.165 0.7 4.165 0.45 0.475 0.45 0.475 1.17 0.245 1.17 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.245 3.28 0.475 3.28 0.475 3.86 8.585 3.86 8.585 3.28 8.815 3.28 8.815 4.09 0.245 4.09  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__aoi211_2
