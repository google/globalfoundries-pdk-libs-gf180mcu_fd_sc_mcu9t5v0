# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__invz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__invz_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 20.72 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.27 1.77 1.555 1.77 1.555 2.71 1.27 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER METAL1 ;
        POLYGON 5.165 2.33 5.45 2.33 5.45 3.27 5.165 3.27  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.6696 ;
    PORT
      LAYER METAL1 ;
        POLYGON 12.215 2.925 17.195 2.925 17.535 2.925 18.315 2.925 18.315 1.595 12.165 1.595 12.165 0.68 12.395 0.68 12.395 1.21 14.405 1.21 14.405 0.68 14.635 0.68 14.635 1.215 16.645 1.215 16.645 0.68 16.875 0.68 16.875 1.21 18.885 1.21 18.885 0.68 19.115 0.68 19.115 1.595 18.805 1.595 18.805 4.195 18.335 4.195 18.335 3.155 17.535 3.155 17.195 3.155 16.525 3.155 16.525 4.195 16.295 4.195 16.295 3.155 14.485 3.155 14.485 4.19 14.255 4.19 14.255 3.155 12.455 3.155 12.455 4.19 12.215 4.19  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.905 4.59 1.905 3.42 2.135 3.42 2.135 4.59 4.675 4.59 4.675 4.35 4.905 4.35 4.905 4.59 6.715 4.59 6.715 4.35 6.945 4.35 6.945 4.59 8.755 4.59 8.755 3.38 8.985 3.38 8.985 4.59 10.995 4.59 10.995 3.88 11.225 3.88 11.225 4.59 13.235 4.59 13.235 3.385 13.465 3.385 13.465 4.59 15.275 4.59 15.275 3.385 15.505 3.385 15.505 4.59 17.195 4.59 17.315 4.59 17.315 3.385 17.535 3.385 17.545 3.385 17.545 4.59 19.355 4.59 19.355 3.38 19.585 3.38 19.585 4.59 20.72 4.59 20.72 5.49 17.535 5.49 17.195 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 20.72 -0.45 20.72 0.45 20.235 0.45 20.235 1.49 20.005 1.49 20.005 0.45 17.995 0.45 17.995 0.98 17.765 0.98 17.765 0.45 15.755 0.45 15.755 0.98 15.525 0.98 15.525 0.45 13.515 0.45 13.515 0.98 13.285 0.98 13.285 0.45 11.275 0.45 11.275 1.49 11.045 1.49 11.045 0.45 9.035 0.45 9.035 1.49 8.805 1.49 8.805 0.45 6.85 0.45 6.85 0.635 6.51 0.635 6.51 0.45 4.61 0.45 4.61 0.635 4.27 0.635 4.27 0.45 1.595 0.45 1.595 1.02 1.365 1.02 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.885 2.94 2.63 2.94 2.63 2.11 1.805 2.11 1.805 1.49 0.245 1.49 0.245 0.68 0.475 0.68 0.475 1.26 2.035 1.26 2.035 1.88 2.86 1.88 2.86 2.425 3.65 2.425 3.65 3.15 2.725 3.15 2.725 3.17 1.115 3.17 1.115 4.19 0.885 4.19  ;
        POLYGON 5.695 2.48 7.155 2.48 7.155 1.595 5.39 1.595 5.39 1.365 7.385 1.365 7.385 2.71 5.925 2.71 5.925 3.66 5.695 3.66  ;
        POLYGON 2.925 3.38 3.155 3.38 3.155 3.89 4.405 3.89 4.405 1.595 3.55 1.595 3.55 1.365 4.635 1.365 4.635 3.89 7.735 3.89 7.735 2.405 17.195 2.405 17.195 2.695 10.105 2.695 10.105 4.19 9.875 4.19 9.875 2.695 7.965 2.695 7.965 4.19 7.735 4.19 7.735 4.12 2.925 4.12  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.905 7.63 0.905 7.63 0.855 7.975 0.855 7.975 1.825 9.925 1.825 9.925 0.84 10.155 0.84 10.155 1.825 17.535 1.825 17.535 2.055 7.745 2.055 7.745 1.135 3.32 1.135 3.32 1.825 4.175 1.825 4.175 3.66 3.945 3.66 3.945 2.055 3.09 2.055 3.09 1.49 2.485 1.49  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__invz_8
