# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__nand2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__nand2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.96 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.67 2.47 3.01 2.47 3.01 2.95 5.73 2.95 5.73 2.47 6.07 2.47 6.07 3.21 2.67 3.21  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.458 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.77 1.83 8.11 1.83 8.11 2.15 0.77 2.15  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.8538 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 3.55 7.385 3.55 7.385 3.23 8.34 3.23 8.34 1.105 7.94 1.105 7.94 1.1 2.275 1.1 2.275 0.87 8.145 0.87 8.145 0.875 8.57 0.875 8.57 3.46 7.75 3.46 7.75 4.33 7.37 4.33 7.37 3.78 5.575 3.78 5.575 4.36 5.345 4.36 5.345 3.78 3.535 3.78 3.535 4.36 3.305 4.36 3.305 3.78 1.495 3.78 1.495 4.36 1.265 4.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.69 0.475 3.69 0.475 4.59 2.285 4.59 2.285 4.16 2.515 4.16 2.515 4.59 4.325 4.59 4.325 4.16 4.555 4.16 4.555 4.59 6.365 4.59 6.365 4.16 6.595 4.16 6.595 4.59 8.405 4.59 8.405 3.69 8.635 3.69 8.635 4.59 8.96 4.59 8.96 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.96 -0.45 8.96 0.45 8.69 0.45 8.69 0.64 8.35 0.64 8.35 0.45 4.575 0.45 4.575 0.64 4.235 0.64 4.235 0.45 0.555 0.45 0.555 1.165 0.325 1.165 0.325 0.45 0 0.45  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu9t5v0__nand2_4
