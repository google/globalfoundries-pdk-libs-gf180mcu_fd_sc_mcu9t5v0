* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__xnor2_2 A1 A2 ZN VDD VNW VPW VSS
*.PININFO A1:I A2:I ZN:O VDD:P VNW:P VPW:P VSS:G
*.EQN ZN=!(!((A1 * A2) + !(A1 + A2)))
M_i_8 I A2 VSS VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_9 VSS A1 I VPW nmos_5p0 W=0.660000U L=0.600000U
M_i_4 Z_neg I VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_2 net_0 A1 Z_neg VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_3 VSS A2 net_0 VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_0 ZN Z_neg VSS VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_0_1 VSS Z_neg ZN VPW nmos_5p0 W=1.320000U L=0.600000U
M_i_10 net_2 A2 I VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_11 VDD A1 net_2 VNW pmos_5p0 W=0.915000U L=0.500000U
M_i_7 net_1 I VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_5 Z_neg A1 net_1 VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_6 net_1 A2 Z_neg VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_0 ZN Z_neg VDD VNW pmos_5p0 W=1.830000U L=0.500000U
M_i_1_1 VDD Z_neg ZN VNW pmos_5p0 W=1.830000U L=0.500000U
.ENDS
