# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__bufz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__bufz_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 25.2 BY 5.04 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.384 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.33 1.575 2.33 1.575 2.71 0.71 2.71  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.152 ;
    PORT
      LAYER METAL1 ;
        POLYGON 6.04 1.77 11.05 1.77 11.05 2.15 6.04 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.7344 ;
    PORT
      LAYER METAL1 ;
        POLYGON 12.255 3.365 21.21 3.365 22.08 3.365 22.08 1.6 12.355 1.6 12.355 0.865 23.785 0.865 23.785 1.65 22.685 1.65 22.685 4.175 21.21 4.175 12.255 4.175  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.505 4.59 1.505 3.845 1.735 3.845 1.735 4.59 5.115 4.59 5.115 3.88 5.345 3.88 5.345 4.59 7.155 4.59 7.155 3.88 7.385 3.88 7.385 4.59 9.195 4.59 9.195 3.88 9.425 3.88 9.425 4.59 11.235 4.59 11.235 3.88 11.465 3.88 11.465 4.59 13.22 4.59 13.22 4.405 13.56 4.405 13.56 4.59 15.26 4.59 15.26 4.405 15.6 4.405 15.6 4.59 17.3 4.59 17.3 4.405 17.64 4.405 17.64 4.59 19.34 4.59 19.34 4.405 19.68 4.405 19.68 4.59 21.21 4.59 21.38 4.59 21.38 4.405 21.72 4.405 21.72 4.59 23.475 4.59 23.475 3.88 23.705 3.88 23.705 4.59 25.2 4.59 25.2 5.49 21.21 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 25.2 -0.45 25.2 0.45 24.905 0.45 24.905 1.16 24.675 1.16 24.675 0.45 22.72 0.45 22.72 0.635 22.38 0.635 22.38 0.45 20.48 0.45 20.48 0.635 20.14 0.635 20.14 0.45 18.24 0.45 18.24 0.635 17.9 0.635 17.9 0.45 16 0.45 16 0.635 15.66 0.635 15.66 0.45 13.76 0.45 13.76 0.635 13.42 0.635 13.42 0.45 11.52 0.45 11.52 0.635 11.18 0.635 11.18 0.45 9.28 0.45 9.28 0.635 8.94 0.635 8.94 0.45 7.04 0.45 7.04 0.635 6.7 0.635 6.7 0.45 4.61 0.45 4.61 0.625 4.27 0.625 4.27 0.45 1.595 0.45 1.595 0.695 1.365 0.695 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.485 2.94 1.805 2.94 1.805 1.6 0.19 1.6 0.19 1.37 2.035 1.37 2.035 2.94 3.365 2.94 3.365 2.415 3.595 2.415 3.595 3.17 0.715 3.17 0.715 3.75 0.485 3.75  ;
        POLYGON 2.485 0.68 2.715 0.68 2.715 0.855 5.865 0.855 5.865 0.865 7.875 0.865 7.875 0.68 8.105 0.68 8.105 1.26 10.115 1.26 10.115 0.68 10.345 0.68 10.345 1.26 11.905 1.26 11.905 1.83 21.035 1.83 21.035 2.15 11.675 2.15 11.675 1.49 5.635 1.49 5.635 1.085 3.375 1.085 3.375 1.955 4.175 1.955 4.175 3.215 3.945 3.215 3.945 2.185 3.145 2.185 3.145 1.49 2.485 1.49  ;
        POLYGON 2.925 3.445 4.405 3.445 4.405 1.655 3.605 1.655 3.605 1.315 4.635 1.315 4.635 2.91 11.465 2.91 11.465 2.45 21.21 2.45 21.21 2.79 11.695 2.79 11.695 3.14 10.445 3.14 10.445 3.94 10.215 3.94 10.215 3.36 4.635 3.36 4.635 3.675 3.155 3.675 3.155 4.255 2.925 4.255  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__bufz_12
