# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 17.36 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.854 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.4 1.69 4.325 1.69 4.325 2.235 3.4 2.235  ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.71 2.33 1.865 2.33 1.865 2.71 0.71 2.71  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER METAL1 ;
        POLYGON 15.71 1.37 16.09 1.37 16.09 3.27 15.82 3.27 15.82 1.6 15.71 1.6  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 1.655 4.59 1.655 3.425 1.885 3.425 1.885 4.59 2.325 4.59 3.495 4.59 3.495 3.615 3.725 3.615 3.725 4.59 6.69 4.59 7.925 4.59 7.925 3.145 8.155 3.145 8.155 4.59 9.495 4.59 12.805 4.59 12.805 4.345 13.035 4.345 13.035 4.59 14.8 4.59 14.8 4.345 15.03 4.345 15.03 4.59 16.55 4.59 16.84 4.59 16.84 3.875 17.07 3.875 17.07 4.59 17.36 4.59 17.36 5.49 16.55 5.49 9.495 5.49 6.69 5.49 2.325 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 17.36 -0.45 17.36 0.45 17.115 0.45 17.115 1.165 16.885 1.165 16.885 0.45 14.93 0.45 14.93 0.64 14.59 0.64 14.59 0.45 13.035 0.45 13.035 1.165 12.805 1.165 12.805 0.45 8.155 0.45 8.155 1.19 7.925 1.19 7.925 0.45 3.625 0.45 3.625 1.19 3.395 1.19 3.395 0.45 1.785 0.45 1.785 1.225 1.555 1.225 1.555 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 0.635 2.94 2.095 2.94 2.095 1.74 0.435 1.74 0.435 1.315 0.665 1.315 0.665 1.51 2.325 1.51 2.325 3.17 0.865 3.17 0.865 3.75 0.635 3.75  ;
        POLYGON 4.515 2.975 4.56 2.975 4.56 1.08 4.79 1.08 4.79 3.785 4.515 3.785  ;
        POLYGON 2.675 1.315 2.905 1.315 2.905 2.985 4.185 2.985 4.185 4.13 6.69 4.13 6.69 4.36 3.955 4.36 3.955 3.215 2.675 3.215  ;
        POLYGON 5.965 1.08 6.195 1.08 6.195 2.055 8.595 2.055 8.595 2.395 8.365 2.395 8.365 2.285 6.195 2.285 6.195 3.785 5.965 3.785  ;
        POLYGON 7.485 2.515 7.715 2.515 7.715 2.625 8.945 2.625 8.945 2.055 9.265 2.055 9.265 1.315 9.495 1.315 9.495 2.285 9.175 2.285 9.175 3.785 8.945 3.785 8.945 2.855 7.485 2.855  ;
        POLYGON 6.59 1.595 8.805 1.595 8.805 0.68 11.4 0.68 11.4 2.19 11.55 2.19 11.55 2.42 11.17 2.42 11.17 0.91 9.035 0.91 9.035 1.825 6.59 1.825  ;
        POLYGON 10.385 1.315 10.615 1.315 10.615 2.65 13.19 2.65 13.19 2.47 13.53 2.47 13.53 2.88 10.615 2.88 10.615 3.785 10.385 3.785  ;
        POLYGON 12.31 1.92 13.87 1.92 13.87 1.37 14.21 1.37 14.21 1.83 15.525 1.83 15.525 2.06 14.055 2.06 14.055 3.215 13.825 3.215 13.825 2.15 12.31 2.15  ;
        POLYGON 11.785 3.11 12.015 3.11 12.015 3.69 16.32 3.69 16.32 1.14 13.64 1.14 13.64 1.625 11.63 1.625 11.63 1.37 11.97 1.37 11.97 1.395 13.41 1.395 13.41 0.91 16.55 0.91 16.55 3.92 11.785 3.92  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffnq_2
