# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__fillcap_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__fillcap_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 8.96 BY 5.04 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.97 4.59 1.765 4.59 1.765 3.55 1.995 3.55 1.995 4.59 3.21 4.59 4.005 4.59 4.005 3.55 4.235 3.55 4.235 4.59 5.45 4.59 6.245 4.59 6.245 3.55 6.475 3.55 6.475 4.59 7.69 4.59 8.485 4.59 8.485 3.55 8.715 3.55 8.715 4.59 8.96 4.59 8.96 5.49 8.715 5.49 7.69 5.49 6.475 5.49 5.45 5.49 4.235 5.49 3.21 5.49 1.995 5.49 0.97 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 8.96 -0.45 8.96 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.83 0.97 1.83 0.97 2.06 0.475 2.06 0.475 4.36 0.245 4.36  ;
        POLYGON 1.27 2.47 1.765 2.47 1.765 0.68 1.995 0.68 1.995 2.7 1.27 2.7  ;
        POLYGON 2.485 1.83 3.21 1.83 3.21 2.06 2.715 2.06 2.715 4.36 2.485 4.36  ;
        POLYGON 3.51 2.47 4.005 2.47 4.005 0.68 4.235 0.68 4.235 2.7 3.51 2.7  ;
        POLYGON 4.725 1.83 5.45 1.83 5.45 2.06 4.955 2.06 4.955 4.36 4.725 4.36  ;
        POLYGON 5.75 2.47 6.245 2.47 6.245 0.68 6.475 0.68 6.475 2.7 5.75 2.7  ;
        POLYGON 6.965 1.83 7.69 1.83 7.69 2.06 7.195 2.06 7.195 4.36 6.965 4.36  ;
        POLYGON 7.99 2.47 8.485 2.47 8.485 0.68 8.715 0.68 8.715 2.7 7.99 2.7  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__fillcap_16
