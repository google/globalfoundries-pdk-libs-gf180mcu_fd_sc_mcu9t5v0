* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.SUBCKT gf180mcu_fd_sc_mcu9t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
*.PININFO D:I CLK:I Q:O VDD:P VNW:P VPW:P VSS:G
M_tn3 VSS CLK ncki VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn4 cki ncki VSS VPW nfet_05v0 W=0.790000U L=0.600000U
M_tn5 net5 ncki VSS VPW nfet_05v0 W=0.580000U L=0.600000U
M_tn8 net4 D net5 VPW nfet_05v0 W=0.580000U L=0.600000U
M_tn6 net6 cki net4 VPW nfet_05v0 W=0.580000U L=0.600000U
M_tn7 VSS net0 net6 VPW nfet_05v0 W=0.580000U L=0.600000U
M_tn0 net0 net4 VSS VPW nfet_05v0 W=0.580000U L=0.600000U
M_tn9 net2 cki net0 VPW nfet_05v0 W=0.580000U L=0.600000U
M_tn11 net1 ncki net2 VPW nfet_05v0 W=0.580000U L=0.600000U
M_tn12 VSS net3 net1 VPW nfet_05v0 W=0.580000U L=0.600000U
M_tn10 net3 net2 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_tn1 Q net3 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_tn1_18 Q net3 VSS VPW nfet_05v0 W=1.320000U L=0.600000U
M_tp3 VDD CLK ncki VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp4 cki ncki VDD VNW pfet_05v0 W=1.380000U L=0.500000U
M_tp12 net7 cki VDD VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp11 net4 D net7 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp6 net8 ncki net4 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp5 VDD net0 net8 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp0 net0 net4 VDD VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp7 net2 ncki net0 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp9 net1x cki net2 VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp10 VDD net3 net1x VNW pfet_05v0 W=1.000000U L=0.500000U
M_tp8 net3 net2 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_tp1 Q net3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
M_tp1_16 Q net3 VDD VNW pfet_05v0 W=1.830000U L=0.500000U
.ENDS
