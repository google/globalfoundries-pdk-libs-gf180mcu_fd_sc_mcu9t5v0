# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__xor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__xor2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 6.72 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 1.905 2.87 1.905 2.87 2.33 3.44 2.33 3.885 2.33 3.885 1.85 4.455 1.85 4.455 2.19 4.115 2.19 4.115 2.71 3.44 2.71 2.64 2.71 2.64 2.135 1.94 2.135  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.5605 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.85 1.015 1.85 1.015 2.94 3.44 2.94 4.345 2.94 4.345 2.47 4.83 2.47 4.83 1.905 5.53 1.905 5.53 2.135 5.06 2.135 5.06 2.7 4.575 2.7 4.575 3.17 3.44 3.17 0.71 3.17  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.805 3.04 5.19 3.04 5.19 2.89 5.76 2.89 5.76 1.62 3.785 1.62 3.785 0.81 4.015 0.81 4.015 1.39 5.99 1.39 5.99 3.12 5.45 3.12 5.45 3.27 5.035 3.27 5.035 3.9 4.805 3.9  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 2.435 4.59 2.435 3.4 2.665 3.4 2.665 4.59 3.44 4.59 6.055 4.59 6.72 4.59 6.72 5.49 6.055 5.49 3.44 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 6.72 -0.45 6.72 0.45 6.055 0.45 6.055 1.16 5.825 1.16 5.825 0.45 2.715 0.45 2.715 1.15 2.485 1.15 2.485 0.45 0.475 0.45 0.475 1.15 0.245 1.15 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.25 1.39 1.365 1.39 1.365 0.81 1.595 0.81 1.595 1.39 3.44 1.39 3.44 2.1 3.1 2.1 3.1 1.62 0.48 1.62 0.48 3.4 0.575 3.4 0.575 3.74 0.25 3.74  ;
        POLYGON 3.785 3.4 4.015 3.4 4.015 4.13 5.825 4.13 5.825 3.4 6.055 3.4 6.055 4.36 3.785 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__xor2_1
