# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__buf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__buf_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 7.84 BY 5.04 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.414 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 2.27 1.91 2.27 1.91 2.65 0.63 2.65  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.642 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.605 3.09 4.62 3.09 5.575 3.09 5.575 1.95 3.605 1.95 3.605 0.68 3.865 0.68 3.865 1.72 5.845 1.72 5.845 0.68 6.075 0.68 6.075 4.36 5.745 4.36 5.745 3.32 4.62 3.32 3.835 3.32 3.835 4.36 3.605 4.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 0.245 4.59 0.245 3.55 0.475 3.55 0.475 4.59 2.385 4.59 2.385 3.55 2.615 3.55 2.615 4.59 4.62 4.59 4.625 4.59 4.625 3.55 4.855 3.55 4.855 4.59 6.865 4.59 6.865 3.55 7.095 3.55 7.095 4.59 7.84 4.59 7.84 5.49 4.62 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 7.84 -0.45 7.84 0.45 7.195 0.45 7.195 1.49 6.965 1.49 6.965 0.45 4.955 0.45 4.955 1.49 4.725 1.49 4.725 0.45 2.715 0.45 2.715 1.49 2.485 1.49 2.485 0.45 0.475 0.45 0.475 1.49 0.245 1.49 0.245 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 3.09 2.14 3.09 2.14 1.92 1.365 1.92 1.365 0.68 1.595 0.68 1.595 1.69 2.37 1.69 2.37 2.27 4.62 2.27 4.62 2.5 2.37 2.5 2.37 3.32 1.595 3.32 1.595 4.36 1.365 4.36  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__buf_4
