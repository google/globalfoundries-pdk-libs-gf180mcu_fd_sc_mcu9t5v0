# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__and2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__and2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 5.04 BY 5.04 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.612 ;
    PORT
      LAYER METAL1 ;
        POLYGON 0.15 2.33 0.71 2.33 0.71 1.905 0.97 1.905 0.97 2.715 0.15 2.715  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.612 ;
    PORT
      LAYER METAL1 ;
        POLYGON 1.27 2.33 1.83 2.33 1.83 1.9 2.09 1.9 2.09 2.71 1.27 2.71  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.638 ;
    PORT
      LAYER METAL1 ;
        POLYGON 3.42 0.845 3.77 0.845 3.77 3.685 3.42 3.685  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 4.59 0.26 4.59 0.26 3.685 0.49 3.685 0.49 4.59 2.52 4.59 2.52 3.875 2.75 3.875 2.75 4.59 2.97 4.59 4.56 4.59 4.56 3.875 4.79 3.875 4.79 4.59 5.04 4.59 5.04 5.49 2.97 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER METAL1 ;
        POLYGON 0 -0.45 5.04 -0.45 5.04 0.45 4.77 0.45 4.77 1.165 4.54 1.165 4.54 0.45 2.53 0.45 2.53 1.165 2.3 1.165 2.3 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER METAL1 ;
        POLYGON 1.28 2.94 2.74 2.94 2.74 1.655 0.26 1.655 0.26 0.845 0.49 0.845 0.49 1.425 2.97 1.425 2.97 3.17 1.51 3.17 1.51 3.75 1.28 3.75  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__and2_2
