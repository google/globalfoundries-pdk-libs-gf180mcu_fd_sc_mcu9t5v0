# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu9t5v0__dffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_green_sc9 ;
  SIZE 19.04 BY 5.04 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.96 2.33 3.895 2.33 3.895 2.71 2.96 2.71  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.255 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.59 2.33 14.015 2.33 14.015 2.71 13.59 2.71  ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.164 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 2.265 1.59 2.265 1.59 2.71 0.71 2.71  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6016 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.445 0.845 17.77 0.845 17.77 3.685 17.445 3.685  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 4.59 1.365 4.59 1.365 3.425 1.595 3.425 1.595 4.59 2.09 4.59 3.225 4.59 3.225 3.615 3.455 3.615 3.455 4.59 4.97 4.59 7.305 4.59 7.305 3.615 7.535 3.615 7.535 4.59 8.555 4.59 9.045 4.59 9.045 3.32 9.275 3.32 9.275 4.59 9.77 4.59 10.295 4.59 13.345 4.59 13.345 4.345 13.575 4.345 13.575 4.59 15.155 4.59 15.385 4.59 15.385 3.875 15.615 3.875 15.615 4.59 16.425 4.59 16.425 3.875 16.655 3.875 16.655 4.59 17.05 4.59 18.465 4.59 18.465 3.875 18.695 3.875 18.695 4.59 19.04 4.59 19.04 5.49 17.05 5.49 15.155 5.49 10.295 5.49 9.77 5.49 8.555 5.49 4.97 5.49 2.09 5.49 0 5.49  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.45 19.04 -0.45 19.04 0.45 18.795 0.45 18.795 1.235 18.565 1.235 18.565 0.45 16.555 0.45 16.555 1.235 16.325 1.235 16.325 0.45 13.365 0.45 13.365 1.195 13.135 1.195 13.135 0.45 8.655 0.45 8.655 1.195 8.425 1.195 8.425 0.45 3.435 0.45 3.435 1.195 3.205 1.195 3.205 0.45 1.595 0.45 1.595 1.2 1.365 1.2 1.365 0.45 0 0.45  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.925 0.575 2.925 0.575 2.965 1.86 2.965 1.86 2.035 0.245 2.035 0.245 1.29 0.475 1.29 0.475 1.805 2.09 1.805 2.09 3.195 0.575 3.195 0.575 3.735 0.345 3.735  ;
        POLYGON 4.245 1.195 4.555 1.195 4.555 3.785 4.245 3.785  ;
        POLYGON 2.385 1.29 2.715 1.29 2.715 3.155 3.915 3.155 3.915 4.13 4.97 4.13 4.97 4.36 3.685 4.36 3.685 3.385 2.615 3.385 2.615 3.685 2.385 3.685  ;
        POLYGON 6.285 3.145 8.555 3.145 8.555 3.955 8.325 3.955 8.325 3.375 6.515 3.375 6.515 3.955 6.285 3.955  ;
        POLYGON 5.495 2.685 9.77 2.685 9.77 2.915 5.495 2.915 5.495 3.785 5.265 3.785 5.265 1.185 5.675 1.185 5.675 1.525 5.495 1.525  ;
        POLYGON 6.81 2.225 9.765 2.225 9.765 1.195 9.995 1.195 9.995 2.225 10.295 2.225 10.295 3.96 10.065 3.96 10.065 2.455 6.81 2.455  ;
        POLYGON 5.855 1.71 9.305 1.71 9.305 0.735 11.785 0.735 11.785 2.69 11.815 2.69 11.815 3.03 11.555 3.03 11.555 0.965 10.455 0.965 10.455 1.995 10.225 1.995 10.225 0.965 9.535 0.965 9.535 1.94 5.855 1.94  ;
        POLYGON 12.015 1.195 12.335 1.195 12.335 3.49 12.105 3.49 12.105 1.535 12.015 1.535  ;
        POLYGON 10.895 1.195 11.315 1.195 11.315 3.73 14.925 3.73 14.925 2.415 15.155 2.415 15.155 3.96 10.895 3.96  ;
        POLYGON 12.63 2.745 12.97 2.745 12.97 2.94 14.465 2.94 14.465 1.955 15.555 1.955 15.555 0.725 15.785 0.725 15.785 1.83 17.05 1.83 17.05 2.185 14.695 2.185 14.695 3.17 12.63 3.17  ;
  END
END gf180mcu_fd_sc_mcu9t5v0__dffrnq_2
